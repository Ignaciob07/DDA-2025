module lut_atan #(
    parameter NB_DATA_IN    = 8,
    parameter NB_DATA_OUT   = 16
) (
    output [NB_DATA_OUT - 1 : 0] o_atan      ,
    input  [NB_DATA_IN  - 1 : 0] i_data_i    ,
    input  [NB_DATA_IN  - 1 : 0] i_data_q    ,
    input                        i_clock       ,
    input                        i_rst_n    
);

    localparam NB_LUT   = 16384; // 
    localparam NB_INDEX = (NB_DATA_IN - 1)* 2          ; //

    reg  [NB_INDEX    - 1 : 0] index                 ;
    reg  [NB_DATA_IN  - 1 : 0] data_i                ;
    reg  [NB_DATA_IN  - 1 : 0] data_q                ;
    reg  [NB_DATA_OUT - 1 : 0] r_atan                ;
    reg  [NB_DATA_OUT - 1 : 0] lut [NB_LUT - 1 : 0];

    always @(*) begin
        if(i_data_i[NB_DATA_IN  - 1])                   
            data_i = ~i_data_i + 1;                     
        else                                            
            data_i = i_data_i;                           

        if(i_data_q[NB_DATA_IN  - 1])                   
            data_q = ~i_data_q + 1;                     
        else                                            
            data_q = i_data_q;                           

        index [13-:7] = data_i;        index [6-:7] = data_q;        r_atan = lut[index];                                 
                                                           
    end

    assign o_atan = r_atan;

    always @(posedge i_clock or negedge i_rst_n) begin
        if (!i_rst_n) begin
          lut[0] <= 0;
          lut[1] <= 0;
          lut[2] <= 0;
          lut[3] <= 0;
          lut[4] <= 0;
          lut[5] <= 0;
          lut[6] <= 0;
          lut[7] <= 0;
          lut[8] <= 0;
          lut[9] <= 0;
          lut[10] <= 0;
          lut[11] <= 0;
          lut[12] <= 0;
          lut[13] <= 0;
          lut[14] <= 0;
          lut[15] <= 0;
          lut[16] <= 0;
          lut[17] <= 0;
          lut[18] <= 0;
          lut[19] <= 0;
          lut[20] <= 0;
          lut[21] <= 0;
          lut[22] <= 0;
          lut[23] <= 0;
          lut[24] <= 0;
          lut[25] <= 0;
          lut[26] <= 0;
          lut[27] <= 0;
          lut[28] <= 0;
          lut[29] <= 0;
          lut[30] <= 0;
          lut[31] <= 0;
          lut[32] <= 0;
          lut[33] <= 0;
          lut[34] <= 0;
          lut[35] <= 0;
          lut[36] <= 0;
          lut[37] <= 0;
          lut[38] <= 0;
          lut[39] <= 0;
          lut[40] <= 0;
          lut[41] <= 0;
          lut[42] <= 0;
          lut[43] <= 0;
          lut[44] <= 0;
          lut[45] <= 0;
          lut[46] <= 0;
          lut[47] <= 0;
          lut[48] <= 0;
          lut[49] <= 0;
          lut[50] <= 0;
          lut[51] <= 0;
          lut[52] <= 0;
          lut[53] <= 0;
          lut[54] <= 0;
          lut[55] <= 0;
          lut[56] <= 0;
          lut[57] <= 0;
          lut[58] <= 0;
          lut[59] <= 0;
          lut[60] <= 0;
          lut[61] <= 0;
          lut[62] <= 0;
          lut[63] <= 0;
          lut[64] <= 0;
          lut[65] <= 0;
          lut[66] <= 0;
          lut[67] <= 0;
          lut[68] <= 0;
          lut[69] <= 0;
          lut[70] <= 0;
          lut[71] <= 0;
          lut[72] <= 0;
          lut[73] <= 0;
          lut[74] <= 0;
          lut[75] <= 0;
          lut[76] <= 0;
          lut[77] <= 0;
          lut[78] <= 0;
          lut[79] <= 0;
          lut[80] <= 0;
          lut[81] <= 0;
          lut[82] <= 0;
          lut[83] <= 0;
          lut[84] <= 0;
          lut[85] <= 0;
          lut[86] <= 0;
          lut[87] <= 0;
          lut[88] <= 0;
          lut[89] <= 0;
          lut[90] <= 0;
          lut[91] <= 0;
          lut[92] <= 0;
          lut[93] <= 0;
          lut[94] <= 0;
          lut[95] <= 0;
          lut[96] <= 0;
          lut[97] <= 0;
          lut[98] <= 0;
          lut[99] <= 0;
          lut[100] <= 0;
          lut[101] <= 0;
          lut[102] <= 0;
          lut[103] <= 0;
          lut[104] <= 0;
          lut[105] <= 0;
          lut[106] <= 0;
          lut[107] <= 0;
          lut[108] <= 0;
          lut[109] <= 0;
          lut[110] <= 0;
          lut[111] <= 0;
          lut[112] <= 0;
          lut[113] <= 0;
          lut[114] <= 0;
          lut[115] <= 0;
          lut[116] <= 0;
          lut[117] <= 0;
          lut[118] <= 0;
          lut[119] <= 0;
          lut[120] <= 0;
          lut[121] <= 0;
          lut[122] <= 0;
          lut[123] <= 0;
          lut[124] <= 0;
          lut[125] <= 0;
          lut[126] <= 0;
          lut[127] <= 0;
          lut[128] <= 0;
          lut[129] <= 16'd12868;
          lut[130] <= 16'd18140;
          lut[131] <= 16'd20464;
          lut[132] <= 16'd21722;
          lut[133] <= 16'd22502;
          lut[134] <= 16'd23030;
          lut[135] <= 16'd23411;
          lut[136] <= 16'd23698;
          lut[137] <= 16'd23923;
          lut[138] <= 16'd24103;
          lut[139] <= 16'd24251;
          lut[140] <= 16'd24374;
          lut[141] <= 16'd24478;
          lut[142] <= 16'd24568;
          lut[143] <= 16'd24645;
          lut[144] <= 16'd24713;
          lut[145] <= 16'd24773;
          lut[146] <= 16'd24827;
          lut[147] <= 16'd24874;
          lut[148] <= 16'd24917;
          lut[149] <= 16'd24956;
          lut[150] <= 16'd24992;
          lut[151] <= 16'd25024;
          lut[152] <= 16'd25054;
          lut[153] <= 16'd25081;
          lut[154] <= 16'd25106;
          lut[155] <= 16'd25129;
          lut[156] <= 16'd25151;
          lut[157] <= 16'd25171;
          lut[158] <= 16'd25190;
          lut[159] <= 16'd25208;
          lut[160] <= 16'd25224;
          lut[161] <= 16'd25240;
          lut[162] <= 16'd25254;
          lut[163] <= 16'd25268;
          lut[164] <= 16'd25281;
          lut[165] <= 16'd25293;
          lut[166] <= 16'd25305;
          lut[167] <= 16'd25316;
          lut[168] <= 16'd25326;
          lut[169] <= 16'd25336;
          lut[170] <= 16'd25346;
          lut[171] <= 16'd25355;
          lut[172] <= 16'd25364;
          lut[173] <= 16'd25372;
          lut[174] <= 16'd25380;
          lut[175] <= 16'd25387;
          lut[176] <= 16'd25395;
          lut[177] <= 16'd25402;
          lut[178] <= 16'd25408;
          lut[179] <= 16'd25415;
          lut[180] <= 16'd25421;
          lut[181] <= 16'd25427;
          lut[182] <= 16'd25433;
          lut[183] <= 16'd25438;
          lut[184] <= 16'd25443;
          lut[185] <= 16'd25449;
          lut[186] <= 16'd25453;
          lut[187] <= 16'd25458;
          lut[188] <= 16'd25463;
          lut[189] <= 16'd25467;
          lut[190] <= 16'd25472;
          lut[191] <= 16'd25476;
          lut[192] <= 16'd25480;
          lut[193] <= 16'd25484;
          lut[194] <= 16'd25488;
          lut[195] <= 16'd25491;
          lut[196] <= 16'd25495;
          lut[197] <= 16'd25498;
          lut[198] <= 16'd25502;
          lut[199] <= 16'd25505;
          lut[200] <= 16'd25508;
          lut[201] <= 16'd25512;
          lut[202] <= 16'd25515;
          lut[203] <= 16'd25517;
          lut[204] <= 16'd25520;
          lut[205] <= 16'd25523;
          lut[206] <= 16'd25526;
          lut[207] <= 16'd25529;
          lut[208] <= 16'd25531;
          lut[209] <= 16'd25534;
          lut[210] <= 16'd25536;
          lut[211] <= 16'd25539;
          lut[212] <= 16'd25541;
          lut[213] <= 16'd25543;
          lut[214] <= 16'd25545;
          lut[215] <= 16'd25548;
          lut[216] <= 16'd25550;
          lut[217] <= 16'd25552;
          lut[218] <= 16'd25554;
          lut[219] <= 16'd25556;
          lut[220] <= 16'd25558;
          lut[221] <= 16'd25560;
          lut[222] <= 16'd25562;
          lut[223] <= 16'd25563;
          lut[224] <= 16'd25565;
          lut[225] <= 16'd25567;
          lut[226] <= 16'd25569;
          lut[227] <= 16'd25570;
          lut[228] <= 16'd25572;
          lut[229] <= 16'd25574;
          lut[230] <= 16'd25575;
          lut[231] <= 16'd25577;
          lut[232] <= 16'd25578;
          lut[233] <= 16'd25580;
          lut[234] <= 16'd25581;
          lut[235] <= 16'd25583;
          lut[236] <= 16'd25584;
          lut[237] <= 16'd25586;
          lut[238] <= 16'd25587;
          lut[239] <= 16'd25588;
          lut[240] <= 16'd25590;
          lut[241] <= 16'd25591;
          lut[242] <= 16'd25592;
          lut[243] <= 16'd25593;
          lut[244] <= 16'd25595;
          lut[245] <= 16'd25596;
          lut[246] <= 16'd25597;
          lut[247] <= 16'd25598;
          lut[248] <= 16'd25599;
          lut[249] <= 16'd25601;
          lut[250] <= 16'd25602;
          lut[251] <= 16'd25603;
          lut[252] <= 16'd25604;
          lut[253] <= 16'd25605;
          lut[254] <= 16'd25606;
          lut[255] <= 16'd25607;
          lut[256] <= 0;
          lut[257] <= 16'd7596;
          lut[258] <= 16'd12868;
          lut[259] <= 16'd16102;
          lut[260] <= 16'd18140;
          lut[261] <= 16'd19502;
          lut[262] <= 16'd20464;
          lut[263] <= 16'd21176;
          lut[264] <= 16'd21722;
          lut[265] <= 16'd22153;
          lut[266] <= 16'd22502;
          lut[267] <= 16'd22789;
          lut[268] <= 16'd23030;
          lut[269] <= 16'd23235;
          lut[270] <= 16'd23411;
          lut[271] <= 16'd23564;
          lut[272] <= 16'd23698;
          lut[273] <= 16'd23817;
          lut[274] <= 16'd23923;
          lut[275] <= 16'd24018;
          lut[276] <= 16'd24103;
          lut[277] <= 16'd24180;
          lut[278] <= 16'd24251;
          lut[279] <= 16'd24315;
          lut[280] <= 16'd24374;
          lut[281] <= 16'd24428;
          lut[282] <= 16'd24478;
          lut[283] <= 16'd24525;
          lut[284] <= 16'd24568;
          lut[285] <= 16'd24608;
          lut[286] <= 16'd24645;
          lut[287] <= 16'd24680;
          lut[288] <= 16'd24713;
          lut[289] <= 16'd24744;
          lut[290] <= 16'd24773;
          lut[291] <= 16'd24801;
          lut[292] <= 16'd24827;
          lut[293] <= 16'd24851;
          lut[294] <= 16'd24874;
          lut[295] <= 16'd24896;
          lut[296] <= 16'd24917;
          lut[297] <= 16'd24937;
          lut[298] <= 16'd24956;
          lut[299] <= 16'd24974;
          lut[300] <= 16'd24992;
          lut[301] <= 16'd25008;
          lut[302] <= 16'd25024;
          lut[303] <= 16'd25039;
          lut[304] <= 16'd25054;
          lut[305] <= 16'd25068;
          lut[306] <= 16'd25081;
          lut[307] <= 16'd25094;
          lut[308] <= 16'd25106;
          lut[309] <= 16'd25118;
          lut[310] <= 16'd25129;
          lut[311] <= 16'd25140;
          lut[312] <= 16'd25151;
          lut[313] <= 16'd25161;
          lut[314] <= 16'd25171;
          lut[315] <= 16'd25181;
          lut[316] <= 16'd25190;
          lut[317] <= 16'd25199;
          lut[318] <= 16'd25208;
          lut[319] <= 16'd25216;
          lut[320] <= 16'd25224;
          lut[321] <= 16'd25232;
          lut[322] <= 16'd25240;
          lut[323] <= 16'd25247;
          lut[324] <= 16'd25254;
          lut[325] <= 16'd25261;
          lut[326] <= 16'd25268;
          lut[327] <= 16'd25275;
          lut[328] <= 16'd25281;
          lut[329] <= 16'd25287;
          lut[330] <= 16'd25293;
          lut[331] <= 16'd25299;
          lut[332] <= 16'd25305;
          lut[333] <= 16'd25310;
          lut[334] <= 16'd25316;
          lut[335] <= 16'd25321;
          lut[336] <= 16'd25326;
          lut[337] <= 16'd25331;
          lut[338] <= 16'd25336;
          lut[339] <= 16'd25341;
          lut[340] <= 16'd25346;
          lut[341] <= 16'd25350;
          lut[342] <= 16'd25355;
          lut[343] <= 16'd25359;
          lut[344] <= 16'd25364;
          lut[345] <= 16'd25368;
          lut[346] <= 16'd25372;
          lut[347] <= 16'd25376;
          lut[348] <= 16'd25380;
          lut[349] <= 16'd25384;
          lut[350] <= 16'd25387;
          lut[351] <= 16'd25391;
          lut[352] <= 16'd25395;
          lut[353] <= 16'd25398;
          lut[354] <= 16'd25402;
          lut[355] <= 16'd25405;
          lut[356] <= 16'd25408;
          lut[357] <= 16'd25412;
          lut[358] <= 16'd25415;
          lut[359] <= 16'd25418;
          lut[360] <= 16'd25421;
          lut[361] <= 16'd25424;
          lut[362] <= 16'd25427;
          lut[363] <= 16'd25430;
          lut[364] <= 16'd25433;
          lut[365] <= 16'd25435;
          lut[366] <= 16'd25438;
          lut[367] <= 16'd25441;
          lut[368] <= 16'd25443;
          lut[369] <= 16'd25446;
          lut[370] <= 16'd25449;
          lut[371] <= 16'd25451;
          lut[372] <= 16'd25453;
          lut[373] <= 16'd25456;
          lut[374] <= 16'd25458;
          lut[375] <= 16'd25461;
          lut[376] <= 16'd25463;
          lut[377] <= 16'd25465;
          lut[378] <= 16'd25467;
          lut[379] <= 16'd25470;
          lut[380] <= 16'd25472;
          lut[381] <= 16'd25474;
          lut[382] <= 16'd25476;
          lut[383] <= 16'd25478;
          lut[384] <= 0;
          lut[385] <= 16'd5272;
          lut[386] <= 16'd9634;
          lut[387] <= 16'd12868;
          lut[388] <= 16'd15193;
          lut[389] <= 16'd16882;
          lut[390] <= 16'd18140;
          lut[391] <= 16'd19102;
          lut[392] <= 16'd19858;
          lut[393] <= 16'd20464;
          lut[394] <= 16'd20961;
          lut[395] <= 16'd21374;
          lut[396] <= 16'd21722;
          lut[397] <= 16'd22020;
          lut[398] <= 16'd22277;
          lut[399] <= 16'd22502;
          lut[400] <= 16'd22699;
          lut[401] <= 16'd22874;
          lut[402] <= 16'd23030;
          lut[403] <= 16'd23170;
          lut[404] <= 16'd23297;
          lut[405] <= 16'd23411;
          lut[406] <= 16'd23515;
          lut[407] <= 16'd23611;
          lut[408] <= 16'd23698;
          lut[409] <= 16'd23779;
          lut[410] <= 16'd23854;
          lut[411] <= 16'd23923;
          lut[412] <= 16'd23987;
          lut[413] <= 16'd24047;
          lut[414] <= 16'd24103;
          lut[415] <= 16'd24155;
          lut[416] <= 16'd24204;
          lut[417] <= 16'd24251;
          lut[418] <= 16'd24294;
          lut[419] <= 16'd24335;
          lut[420] <= 16'd24374;
          lut[421] <= 16'd24410;
          lut[422] <= 16'd24445;
          lut[423] <= 16'd24478;
          lut[424] <= 16'd24509;
          lut[425] <= 16'd24539;
          lut[426] <= 16'd24568;
          lut[427] <= 16'd24595;
          lut[428] <= 16'd24621;
          lut[429] <= 16'd24645;
          lut[430] <= 16'd24669;
          lut[431] <= 16'd24692;
          lut[432] <= 16'd24713;
          lut[433] <= 16'd24734;
          lut[434] <= 16'd24754;
          lut[435] <= 16'd24773;
          lut[436] <= 16'd24792;
          lut[437] <= 16'd24810;
          lut[438] <= 16'd24827;
          lut[439] <= 16'd24843;
          lut[440] <= 16'd24859;
          lut[441] <= 16'd24874;
          lut[442] <= 16'd24889;
          lut[443] <= 16'd24904;
          lut[444] <= 16'd24917;
          lut[445] <= 16'd24931;
          lut[446] <= 16'd24944;
          lut[447] <= 16'd24956;
          lut[448] <= 16'd24968;
          lut[449] <= 16'd24980;
          lut[450] <= 16'd24992;
          lut[451] <= 16'd25003;
          lut[452] <= 16'd25014;
          lut[453] <= 16'd25024;
          lut[454] <= 16'd25034;
          lut[455] <= 16'd25044;
          lut[456] <= 16'd25054;
          lut[457] <= 16'd25063;
          lut[458] <= 16'd25072;
          lut[459] <= 16'd25081;
          lut[460] <= 16'd25090;
          lut[461] <= 16'd25098;
          lut[462] <= 16'd25106;
          lut[463] <= 16'd25114;
          lut[464] <= 16'd25122;
          lut[465] <= 16'd25129;
          lut[466] <= 16'd25137;
          lut[467] <= 16'd25144;
          lut[468] <= 16'd25151;
          lut[469] <= 16'd25158;
          lut[470] <= 16'd25165;
          lut[471] <= 16'd25171;
          lut[472] <= 16'd25178;
          lut[473] <= 16'd25184;
          lut[474] <= 16'd25190;
          lut[475] <= 16'd25196;
          lut[476] <= 16'd25202;
          lut[477] <= 16'd25208;
          lut[478] <= 16'd25213;
          lut[479] <= 16'd25219;
          lut[480] <= 16'd25224;
          lut[481] <= 16'd25229;
          lut[482] <= 16'd25235;
          lut[483] <= 16'd25240;
          lut[484] <= 16'd25245;
          lut[485] <= 16'd25249;
          lut[486] <= 16'd25254;
          lut[487] <= 16'd25259;
          lut[488] <= 16'd25263;
          lut[489] <= 16'd25268;
          lut[490] <= 16'd25272;
          lut[491] <= 16'd25277;
          lut[492] <= 16'd25281;
          lut[493] <= 16'd25285;
          lut[494] <= 16'd25289;
          lut[495] <= 16'd25293;
          lut[496] <= 16'd25297;
          lut[497] <= 16'd25301;
          lut[498] <= 16'd25305;
          lut[499] <= 16'd25309;
          lut[500] <= 16'd25312;
          lut[501] <= 16'd25316;
          lut[502] <= 16'd25319;
          lut[503] <= 16'd25323;
          lut[504] <= 16'd25326;
          lut[505] <= 16'd25330;
          lut[506] <= 16'd25333;
          lut[507] <= 16'd25336;
          lut[508] <= 16'd25340;
          lut[509] <= 16'd25343;
          lut[510] <= 16'd25346;
          lut[511] <= 16'd25349;
          lut[512] <= 0;
          lut[513] <= 16'd4014;
          lut[514] <= 16'd7596;
          lut[515] <= 16'd10543;
          lut[516] <= 16'd12868;
          lut[517] <= 16'd14681;
          lut[518] <= 16'd16102;
          lut[519] <= 16'd17230;
          lut[520] <= 16'd18140;
          lut[521] <= 16'd18884;
          lut[522] <= 16'd19502;
          lut[523] <= 16'd20022;
          lut[524] <= 16'd20464;
          lut[525] <= 16'd20845;
          lut[526] <= 16'd21176;
          lut[527] <= 16'd21466;
          lut[528] <= 16'd21722;
          lut[529] <= 16'd21950;
          lut[530] <= 16'd22153;
          lut[531] <= 16'd22336;
          lut[532] <= 16'd22502;
          lut[533] <= 16'd22652;
          lut[534] <= 16'd22789;
          lut[535] <= 16'd22915;
          lut[536] <= 16'd23030;
          lut[537] <= 16'd23137;
          lut[538] <= 16'd23235;
          lut[539] <= 16'd23326;
          lut[540] <= 16'd23411;
          lut[541] <= 16'd23490;
          lut[542] <= 16'd23564;
          lut[543] <= 16'd23633;
          lut[544] <= 16'd23698;
          lut[545] <= 16'd23760;
          lut[546] <= 16'd23817;
          lut[547] <= 16'd23872;
          lut[548] <= 16'd23923;
          lut[549] <= 16'd23972;
          lut[550] <= 16'd24018;
          lut[551] <= 16'd24061;
          lut[552] <= 16'd24103;
          lut[553] <= 16'd24143;
          lut[554] <= 16'd24180;
          lut[555] <= 16'd24216;
          lut[556] <= 16'd24251;
          lut[557] <= 16'd24283;
          lut[558] <= 16'd24315;
          lut[559] <= 16'd24345;
          lut[560] <= 16'd24374;
          lut[561] <= 16'd24401;
          lut[562] <= 16'd24428;
          lut[563] <= 16'd24454;
          lut[564] <= 16'd24478;
          lut[565] <= 16'd24502;
          lut[566] <= 16'd24525;
          lut[567] <= 16'd24546;
          lut[568] <= 16'd24568;
          lut[569] <= 16'd24588;
          lut[570] <= 16'd24608;
          lut[571] <= 16'd24627;
          lut[572] <= 16'd24645;
          lut[573] <= 16'd24663;
          lut[574] <= 16'd24680;
          lut[575] <= 16'd24697;
          lut[576] <= 16'd24713;
          lut[577] <= 16'd24729;
          lut[578] <= 16'd24744;
          lut[579] <= 16'd24759;
          lut[580] <= 16'd24773;
          lut[581] <= 16'd24787;
          lut[582] <= 16'd24801;
          lut[583] <= 16'd24814;
          lut[584] <= 16'd24827;
          lut[585] <= 16'd24839;
          lut[586] <= 16'd24851;
          lut[587] <= 16'd24863;
          lut[588] <= 16'd24874;
          lut[589] <= 16'd24886;
          lut[590] <= 16'd24896;
          lut[591] <= 16'd24907;
          lut[592] <= 16'd24917;
          lut[593] <= 16'd24927;
          lut[594] <= 16'd24937;
          lut[595] <= 16'd24947;
          lut[596] <= 16'd24956;
          lut[597] <= 16'd24965;
          lut[598] <= 16'd24974;
          lut[599] <= 16'd24983;
          lut[600] <= 16'd24992;
          lut[601] <= 16'd25000;
          lut[602] <= 16'd25008;
          lut[603] <= 16'd25016;
          lut[604] <= 16'd25024;
          lut[605] <= 16'd25032;
          lut[606] <= 16'd25039;
          lut[607] <= 16'd25046;
          lut[608] <= 16'd25054;
          lut[609] <= 16'd25061;
          lut[610] <= 16'd25068;
          lut[611] <= 16'd25074;
          lut[612] <= 16'd25081;
          lut[613] <= 16'd25087;
          lut[614] <= 16'd25094;
          lut[615] <= 16'd25100;
          lut[616] <= 16'd25106;
          lut[617] <= 16'd25112;
          lut[618] <= 16'd25118;
          lut[619] <= 16'd25124;
          lut[620] <= 16'd25129;
          lut[621] <= 16'd25135;
          lut[622] <= 16'd25140;
          lut[623] <= 16'd25146;
          lut[624] <= 16'd25151;
          lut[625] <= 16'd25156;
          lut[626] <= 16'd25161;
          lut[627] <= 16'd25166;
          lut[628] <= 16'd25171;
          lut[629] <= 16'd25176;
          lut[630] <= 16'd25181;
          lut[631] <= 16'd25185;
          lut[632] <= 16'd25190;
          lut[633] <= 16'd25195;
          lut[634] <= 16'd25199;
          lut[635] <= 16'd25203;
          lut[636] <= 16'd25208;
          lut[637] <= 16'd25212;
          lut[638] <= 16'd25216;
          lut[639] <= 16'd25220;
          lut[640] <= 0;
          lut[641] <= 16'd3234;
          lut[642] <= 16'd6234;
          lut[643] <= 16'd8854;
          lut[644] <= 16'd11055;
          lut[645] <= 16'd12868;
          lut[646] <= 16'd14353;
          lut[647] <= 16'd15574;
          lut[648] <= 16'd16584;
          lut[649] <= 16'd17428;
          lut[650] <= 16'd18140;
          lut[651] <= 16'd18746;
          lut[652] <= 16'd19268;
          lut[653] <= 16'd19720;
          lut[654] <= 16'd20116;
          lut[655] <= 16'd20464;
          lut[656] <= 16'd20773;
          lut[657] <= 16'd21049;
          lut[658] <= 16'd21297;
          lut[659] <= 16'd21520;
          lut[660] <= 16'd21722;
          lut[661] <= 16'd21906;
          lut[662] <= 16'd22074;
          lut[663] <= 16'd22229;
          lut[664] <= 16'd22371;
          lut[665] <= 16'd22502;
          lut[666] <= 16'd22623;
          lut[667] <= 16'd22736;
          lut[668] <= 16'd22841;
          lut[669] <= 16'd22939;
          lut[670] <= 16'd23030;
          lut[671] <= 16'd23116;
          lut[672] <= 16'd23196;
          lut[673] <= 16'd23272;
          lut[674] <= 16'd23344;
          lut[675] <= 16'd23411;
          lut[676] <= 16'd23475;
          lut[677] <= 16'd23535;
          lut[678] <= 16'd23592;
          lut[679] <= 16'd23647;
          lut[680] <= 16'd23698;
          lut[681] <= 16'd23748;
          lut[682] <= 16'd23795;
          lut[683] <= 16'd23839;
          lut[684] <= 16'd23882;
          lut[685] <= 16'd23923;
          lut[686] <= 16'd23962;
          lut[687] <= 16'd23999;
          lut[688] <= 16'd24035;
          lut[689] <= 16'd24070;
          lut[690] <= 16'd24103;
          lut[691] <= 16'd24135;
          lut[692] <= 16'd24165;
          lut[693] <= 16'd24195;
          lut[694] <= 16'd24223;
          lut[695] <= 16'd24251;
          lut[696] <= 16'd24277;
          lut[697] <= 16'd24302;
          lut[698] <= 16'd24327;
          lut[699] <= 16'd24351;
          lut[700] <= 16'd24374;
          lut[701] <= 16'd24396;
          lut[702] <= 16'd24417;
          lut[703] <= 16'd24438;
          lut[704] <= 16'd24459;
          lut[705] <= 16'd24478;
          lut[706] <= 16'd24497;
          lut[707] <= 16'd24516;
          lut[708] <= 16'd24533;
          lut[709] <= 16'd24551;
          lut[710] <= 16'd24568;
          lut[711] <= 16'd24584;
          lut[712] <= 16'd24600;
          lut[713] <= 16'd24615;
          lut[714] <= 16'd24631;
          lut[715] <= 16'd24645;
          lut[716] <= 16'd24660;
          lut[717] <= 16'd24674;
          lut[718] <= 16'd24687;
          lut[719] <= 16'd24700;
          lut[720] <= 16'd24713;
          lut[721] <= 16'd24726;
          lut[722] <= 16'd24738;
          lut[723] <= 16'd24750;
          lut[724] <= 16'd24762;
          lut[725] <= 16'd24773;
          lut[726] <= 16'd24784;
          lut[727] <= 16'd24795;
          lut[728] <= 16'd24806;
          lut[729] <= 16'd24816;
          lut[730] <= 16'd24827;
          lut[731] <= 16'd24837;
          lut[732] <= 16'd24846;
          lut[733] <= 16'd24856;
          lut[734] <= 16'd24865;
          lut[735] <= 16'd24874;
          lut[736] <= 16'd24883;
          lut[737] <= 16'd24892;
          lut[738] <= 16'd24901;
          lut[739] <= 16'd24909;
          lut[740] <= 16'd24917;
          lut[741] <= 16'd24925;
          lut[742] <= 16'd24933;
          lut[743] <= 16'd24941;
          lut[744] <= 16'd24949;
          lut[745] <= 16'd24956;
          lut[746] <= 16'd24964;
          lut[747] <= 16'd24971;
          lut[748] <= 16'd24978;
          lut[749] <= 16'd24985;
          lut[750] <= 16'd24992;
          lut[751] <= 16'd24998;
          lut[752] <= 16'd25005;
          lut[753] <= 16'd25011;
          lut[754] <= 16'd25018;
          lut[755] <= 16'd25024;
          lut[756] <= 16'd25030;
          lut[757] <= 16'd25036;
          lut[758] <= 16'd25042;
          lut[759] <= 16'd25048;
          lut[760] <= 16'd25054;
          lut[761] <= 16'd25059;
          lut[762] <= 16'd25065;
          lut[763] <= 16'd25070;
          lut[764] <= 16'd25076;
          lut[765] <= 16'd25081;
          lut[766] <= 16'd25086;
          lut[767] <= 16'd25091;
          lut[768] <= 0;
          lut[769] <= 16'd2706;
          lut[770] <= 16'd5272;
          lut[771] <= 16'd7596;
          lut[772] <= 16'd9634;
          lut[773] <= 16'd11383;
          lut[774] <= 16'd12868;
          lut[775] <= 16'd14126;
          lut[776] <= 16'd15193;
          lut[777] <= 16'd16102;
          lut[778] <= 16'd16882;
          lut[779] <= 16'd17555;
          lut[780] <= 16'd18140;
          lut[781] <= 16'd18651;
          lut[782] <= 16'd19102;
          lut[783] <= 16'd19502;
          lut[784] <= 16'd19858;
          lut[785] <= 16'd20177;
          lut[786] <= 16'd20464;
          lut[787] <= 16'd20724;
          lut[788] <= 16'd20961;
          lut[789] <= 16'd21176;
          lut[790] <= 16'd21374;
          lut[791] <= 16'd21555;
          lut[792] <= 16'd21722;
          lut[793] <= 16'd21877;
          lut[794] <= 16'd22020;
          lut[795] <= 16'd22153;
          lut[796] <= 16'd22277;
          lut[797] <= 16'd22393;
          lut[798] <= 16'd22502;
          lut[799] <= 16'd22604;
          lut[800] <= 16'd22699;
          lut[801] <= 16'd22789;
          lut[802] <= 16'd22874;
          lut[803] <= 16'd22954;
          lut[804] <= 16'd23030;
          lut[805] <= 16'd23102;
          lut[806] <= 16'd23170;
          lut[807] <= 16'd23235;
          lut[808] <= 16'd23297;
          lut[809] <= 16'd23355;
          lut[810] <= 16'd23411;
          lut[811] <= 16'd23464;
          lut[812] <= 16'd23515;
          lut[813] <= 16'd23564;
          lut[814] <= 16'd23611;
          lut[815] <= 16'd23656;
          lut[816] <= 16'd23698;
          lut[817] <= 16'd23740;
          lut[818] <= 16'd23779;
          lut[819] <= 16'd23817;
          lut[820] <= 16'd23854;
          lut[821] <= 16'd23889;
          lut[822] <= 16'd23923;
          lut[823] <= 16'd23956;
          lut[824] <= 16'd23987;
          lut[825] <= 16'd24018;
          lut[826] <= 16'd24047;
          lut[827] <= 16'd24075;
          lut[828] <= 16'd24103;
          lut[829] <= 16'd24130;
          lut[830] <= 16'd24155;
          lut[831] <= 16'd24180;
          lut[832] <= 16'd24204;
          lut[833] <= 16'd24228;
          lut[834] <= 16'd24251;
          lut[835] <= 16'd24273;
          lut[836] <= 16'd24294;
          lut[837] <= 16'd24315;
          lut[838] <= 16'd24335;
          lut[839] <= 16'd24355;
          lut[840] <= 16'd24374;
          lut[841] <= 16'd24392;
          lut[842] <= 16'd24410;
          lut[843] <= 16'd24428;
          lut[844] <= 16'd24445;
          lut[845] <= 16'd24462;
          lut[846] <= 16'd24478;
          lut[847] <= 16'd24494;
          lut[848] <= 16'd24509;
          lut[849] <= 16'd24525;
          lut[850] <= 16'd24539;
          lut[851] <= 16'd24554;
          lut[852] <= 16'd24568;
          lut[853] <= 16'd24581;
          lut[854] <= 16'd24595;
          lut[855] <= 16'd24608;
          lut[856] <= 16'd24621;
          lut[857] <= 16'd24633;
          lut[858] <= 16'd24645;
          lut[859] <= 16'd24657;
          lut[860] <= 16'd24669;
          lut[861] <= 16'd24680;
          lut[862] <= 16'd24692;
          lut[863] <= 16'd24703;
          lut[864] <= 16'd24713;
          lut[865] <= 16'd24724;
          lut[866] <= 16'd24734;
          lut[867] <= 16'd24744;
          lut[868] <= 16'd24754;
          lut[869] <= 16'd24764;
          lut[870] <= 16'd24773;
          lut[871] <= 16'd24783;
          lut[872] <= 16'd24792;
          lut[873] <= 16'd24801;
          lut[874] <= 16'd24810;
          lut[875] <= 16'd24818;
          lut[876] <= 16'd24827;
          lut[877] <= 16'd24835;
          lut[878] <= 16'd24843;
          lut[879] <= 16'd24851;
          lut[880] <= 16'd24859;
          lut[881] <= 16'd24867;
          lut[882] <= 16'd24874;
          lut[883] <= 16'd24882;
          lut[884] <= 16'd24889;
          lut[885] <= 16'd24896;
          lut[886] <= 16'd24904;
          lut[887] <= 16'd24911;
          lut[888] <= 16'd24917;
          lut[889] <= 16'd24924;
          lut[890] <= 16'd24931;
          lut[891] <= 16'd24937;
          lut[892] <= 16'd24944;
          lut[893] <= 16'd24950;
          lut[894] <= 16'd24956;
          lut[895] <= 16'd24962;
          lut[896] <= 0;
          lut[897] <= 16'd2325;
          lut[898] <= 16'd4560;
          lut[899] <= 16'd6634;
          lut[900] <= 16'd8506;
          lut[901] <= 16'd10162;
          lut[902] <= 16'd11610;
          lut[903] <= 16'd12868;
          lut[904] <= 16'd13959;
          lut[905] <= 16'd14905;
          lut[906] <= 16'd15730;
          lut[907] <= 16'd16451;
          lut[908] <= 16'd17084;
          lut[909] <= 16'd17643;
          lut[910] <= 16'd18140;
          lut[911] <= 16'd18582;
          lut[912] <= 16'd18979;
          lut[913] <= 16'd19336;
          lut[914] <= 16'd19659;
          lut[915] <= 16'd19953;
          lut[916] <= 16'd20220;
          lut[917] <= 16'd20464;
          lut[918] <= 16'd20689;
          lut[919] <= 16'd20895;
          lut[920] <= 16'd21086;
          lut[921] <= 16'd21263;
          lut[922] <= 16'd21427;
          lut[923] <= 16'd21580;
          lut[924] <= 16'd21722;
          lut[925] <= 16'd21855;
          lut[926] <= 16'd21980;
          lut[927] <= 16'd22097;
          lut[928] <= 16'd22208;
          lut[929] <= 16'd22311;
          lut[930] <= 16'd22409;
          lut[931] <= 16'd22502;
          lut[932] <= 16'd22589;
          lut[933] <= 16'd22672;
          lut[934] <= 16'd22751;
          lut[935] <= 16'd22826;
          lut[936] <= 16'd22897;
          lut[937] <= 16'd22965;
          lut[938] <= 16'd23030;
          lut[939] <= 16'd23092;
          lut[940] <= 16'd23151;
          lut[941] <= 16'd23208;
          lut[942] <= 16'd23262;
          lut[943] <= 16'd23314;
          lut[944] <= 16'd23363;
          lut[945] <= 16'd23411;
          lut[946] <= 16'd23457;
          lut[947] <= 16'd23501;
          lut[948] <= 16'd23544;
          lut[949] <= 16'd23584;
          lut[950] <= 16'd23624;
          lut[951] <= 16'd23662;
          lut[952] <= 16'd23698;
          lut[953] <= 16'd23734;
          lut[954] <= 16'd23768;
          lut[955] <= 16'd23801;
          lut[956] <= 16'd23833;
          lut[957] <= 16'd23864;
          lut[958] <= 16'd23894;
          lut[959] <= 16'd23923;
          lut[960] <= 16'd23951;
          lut[961] <= 16'd23978;
          lut[962] <= 16'd24005;
          lut[963] <= 16'd24030;
          lut[964] <= 16'd24055;
          lut[965] <= 16'd24079;
          lut[966] <= 16'd24103;
          lut[967] <= 16'd24126;
          lut[968] <= 16'd24148;
          lut[969] <= 16'd24170;
          lut[970] <= 16'd24191;
          lut[971] <= 16'd24211;
          lut[972] <= 16'd24231;
          lut[973] <= 16'd24251;
          lut[974] <= 16'd24269;
          lut[975] <= 16'd24288;
          lut[976] <= 16'd24306;
          lut[977] <= 16'd24324;
          lut[978] <= 16'd24341;
          lut[979] <= 16'd24357;
          lut[980] <= 16'd24374;
          lut[981] <= 16'd24390;
          lut[982] <= 16'd24405;
          lut[983] <= 16'd24421;
          lut[984] <= 16'd24435;
          lut[985] <= 16'd24450;
          lut[986] <= 16'd24464;
          lut[987] <= 16'd24478;
          lut[988] <= 16'd24492;
          lut[989] <= 16'd24505;
          lut[990] <= 16'd24518;
          lut[991] <= 16'd24531;
          lut[992] <= 16'd24543;
          lut[993] <= 16'd24556;
          lut[994] <= 16'd24568;
          lut[995] <= 16'd24579;
          lut[996] <= 16'd24591;
          lut[997] <= 16'd24602;
          lut[998] <= 16'd24613;
          lut[999] <= 16'd24624;
          lut[1000] <= 16'd24635;
          lut[1001] <= 16'd24645;
          lut[1002] <= 16'd24656;
          lut[1003] <= 16'd24666;
          lut[1004] <= 16'd24675;
          lut[1005] <= 16'd24685;
          lut[1006] <= 16'd24695;
          lut[1007] <= 16'd24704;
          lut[1008] <= 16'd24713;
          lut[1009] <= 16'd24722;
          lut[1010] <= 16'd24731;
          lut[1011] <= 16'd24740;
          lut[1012] <= 16'd24748;
          lut[1013] <= 16'd24757;
          lut[1014] <= 16'd24765;
          lut[1015] <= 16'd24773;
          lut[1016] <= 16'd24781;
          lut[1017] <= 16'd24789;
          lut[1018] <= 16'd24797;
          lut[1019] <= 16'd24805;
          lut[1020] <= 16'd24812;
          lut[1021] <= 16'd24819;
          lut[1022] <= 16'd24827;
          lut[1023] <= 16'd24834;
          lut[1024] <= 0;
          lut[1025] <= 16'd2037;
          lut[1026] <= 16'd4014;
          lut[1027] <= 16'd5878;
          lut[1028] <= 16'd7596;
          lut[1029] <= 16'd9152;
          lut[1030] <= 16'd10543;
          lut[1031] <= 16'd11777;
          lut[1032] <= 16'd12868;
          lut[1033] <= 16'd13831;
          lut[1034] <= 16'd14681;
          lut[1035] <= 16'd15434;
          lut[1036] <= 16'd16102;
          lut[1037] <= 16'd16698;
          lut[1038] <= 16'd17230;
          lut[1039] <= 16'd17708;
          lut[1040] <= 16'd18140;
          lut[1041] <= 16'd18530;
          lut[1042] <= 16'd18884;
          lut[1043] <= 16'd19207;
          lut[1044] <= 16'd19502;
          lut[1045] <= 16'd19772;
          lut[1046] <= 16'd20022;
          lut[1047] <= 16'd20252;
          lut[1048] <= 16'd20464;
          lut[1049] <= 16'd20662;
          lut[1050] <= 16'd20845;
          lut[1051] <= 16'd21016;
          lut[1052] <= 16'd21176;
          lut[1053] <= 16'd21326;
          lut[1054] <= 16'd21466;
          lut[1055] <= 16'd21598;
          lut[1056] <= 16'd21722;
          lut[1057] <= 16'd21839;
          lut[1058] <= 16'd21950;
          lut[1059] <= 16'd22054;
          lut[1060] <= 16'd22153;
          lut[1061] <= 16'd22247;
          lut[1062] <= 16'd22336;
          lut[1063] <= 16'd22421;
          lut[1064] <= 16'd22502;
          lut[1065] <= 16'd22579;
          lut[1066] <= 16'd22652;
          lut[1067] <= 16'd22722;
          lut[1068] <= 16'd22789;
          lut[1069] <= 16'd22853;
          lut[1070] <= 16'd22915;
          lut[1071] <= 16'd22974;
          lut[1072] <= 16'd23030;
          lut[1073] <= 16'd23084;
          lut[1074] <= 16'd23137;
          lut[1075] <= 16'd23187;
          lut[1076] <= 16'd23235;
          lut[1077] <= 16'd23281;
          lut[1078] <= 16'd23326;
          lut[1079] <= 16'd23369;
          lut[1080] <= 16'd23411;
          lut[1081] <= 16'd23451;
          lut[1082] <= 16'd23490;
          lut[1083] <= 16'd23528;
          lut[1084] <= 16'd23564;
          lut[1085] <= 16'd23599;
          lut[1086] <= 16'd23633;
          lut[1087] <= 16'd23666;
          lut[1088] <= 16'd23698;
          lut[1089] <= 16'd23730;
          lut[1090] <= 16'd23760;
          lut[1091] <= 16'd23789;
          lut[1092] <= 16'd23817;
          lut[1093] <= 16'd23845;
          lut[1094] <= 16'd23872;
          lut[1095] <= 16'd23898;
          lut[1096] <= 16'd23923;
          lut[1097] <= 16'd23948;
          lut[1098] <= 16'd23972;
          lut[1099] <= 16'd23995;
          lut[1100] <= 16'd24018;
          lut[1101] <= 16'd24040;
          lut[1102] <= 16'd24061;
          lut[1103] <= 16'd24082;
          lut[1104] <= 16'd24103;
          lut[1105] <= 16'd24123;
          lut[1106] <= 16'd24143;
          lut[1107] <= 16'd24162;
          lut[1108] <= 16'd24180;
          lut[1109] <= 16'd24198;
          lut[1110] <= 16'd24216;
          lut[1111] <= 16'd24234;
          lut[1112] <= 16'd24251;
          lut[1113] <= 16'd24267;
          lut[1114] <= 16'd24283;
          lut[1115] <= 16'd24299;
          lut[1116] <= 16'd24315;
          lut[1117] <= 16'd24330;
          lut[1118] <= 16'd24345;
          lut[1119] <= 16'd24359;
          lut[1120] <= 16'd24374;
          lut[1121] <= 16'd24388;
          lut[1122] <= 16'd24401;
          lut[1123] <= 16'd24415;
          lut[1124] <= 16'd24428;
          lut[1125] <= 16'd24441;
          lut[1126] <= 16'd24454;
          lut[1127] <= 16'd24466;
          lut[1128] <= 16'd24478;
          lut[1129] <= 16'd24490;
          lut[1130] <= 16'd24502;
          lut[1131] <= 16'd24513;
          lut[1132] <= 16'd24525;
          lut[1133] <= 16'd24536;
          lut[1134] <= 16'd24546;
          lut[1135] <= 16'd24557;
          lut[1136] <= 16'd24568;
          lut[1137] <= 16'd24578;
          lut[1138] <= 16'd24588;
          lut[1139] <= 16'd24598;
          lut[1140] <= 16'd24608;
          lut[1141] <= 16'd24617;
          lut[1142] <= 16'd24627;
          lut[1143] <= 16'd24636;
          lut[1144] <= 16'd24645;
          lut[1145] <= 16'd24654;
          lut[1146] <= 16'd24663;
          lut[1147] <= 16'd24672;
          lut[1148] <= 16'd24680;
          lut[1149] <= 16'd24689;
          lut[1150] <= 16'd24697;
          lut[1151] <= 16'd24705;
          lut[1152] <= 0;
          lut[1153] <= 16'd1813;
          lut[1154] <= 16'd3583;
          lut[1155] <= 16'd5272;
          lut[1156] <= 16'd6852;
          lut[1157] <= 16'd8308;
          lut[1158] <= 16'd9634;
          lut[1159] <= 16'd10831;
          lut[1160] <= 16'd11905;
          lut[1161] <= 16'd12868;
          lut[1162] <= 16'd13729;
          lut[1163] <= 16'd14501;
          lut[1164] <= 16'd15193;
          lut[1165] <= 16'd15815;
          lut[1166] <= 16'd16375;
          lut[1167] <= 16'd16882;
          lut[1168] <= 16'd17341;
          lut[1169] <= 16'd17759;
          lut[1170] <= 16'd18140;
          lut[1171] <= 16'd18488;
          lut[1172] <= 16'd18808;
          lut[1173] <= 16'd19102;
          lut[1174] <= 16'd19374;
          lut[1175] <= 16'd19625;
          lut[1176] <= 16'd19858;
          lut[1177] <= 16'd20074;
          lut[1178] <= 16'd20276;
          lut[1179] <= 16'd20464;
          lut[1180] <= 16'd20641;
          lut[1181] <= 16'd20806;
          lut[1182] <= 16'd20961;
          lut[1183] <= 16'd21107;
          lut[1184] <= 16'd21244;
          lut[1185] <= 16'd21374;
          lut[1186] <= 16'd21496;
          lut[1187] <= 16'd21612;
          lut[1188] <= 16'd21722;
          lut[1189] <= 16'd21827;
          lut[1190] <= 16'd21926;
          lut[1191] <= 16'd22020;
          lut[1192] <= 16'd22110;
          lut[1193] <= 16'd22196;
          lut[1194] <= 16'd22277;
          lut[1195] <= 16'd22356;
          lut[1196] <= 16'd22430;
          lut[1197] <= 16'd22502;
          lut[1198] <= 16'd22570;
          lut[1199] <= 16'd22636;
          lut[1200] <= 16'd22699;
          lut[1201] <= 16'd22760;
          lut[1202] <= 16'd22818;
          lut[1203] <= 16'd22874;
          lut[1204] <= 16'd22928;
          lut[1205] <= 16'd22980;
          lut[1206] <= 16'd23030;
          lut[1207] <= 16'd23078;
          lut[1208] <= 16'd23125;
          lut[1209] <= 16'd23170;
          lut[1210] <= 16'd23214;
          lut[1211] <= 16'd23256;
          lut[1212] <= 16'd23297;
          lut[1213] <= 16'd23336;
          lut[1214] <= 16'd23374;
          lut[1215] <= 16'd23411;
          lut[1216] <= 16'd23447;
          lut[1217] <= 16'd23482;
          lut[1218] <= 16'd23515;
          lut[1219] <= 16'd23548;
          lut[1220] <= 16'd23580;
          lut[1221] <= 16'd23611;
          lut[1222] <= 16'd23641;
          lut[1223] <= 16'd23670;
          lut[1224] <= 16'd23698;
          lut[1225] <= 16'd23726;
          lut[1226] <= 16'd23753;
          lut[1227] <= 16'd23779;
          lut[1228] <= 16'd23805;
          lut[1229] <= 16'd23830;
          lut[1230] <= 16'd23854;
          lut[1231] <= 16'd23877;
          lut[1232] <= 16'd23900;
          lut[1233] <= 16'd23923;
          lut[1234] <= 16'd23945;
          lut[1235] <= 16'd23966;
          lut[1236] <= 16'd23987;
          lut[1237] <= 16'd24008;
          lut[1238] <= 16'd24028;
          lut[1239] <= 16'd24047;
          lut[1240] <= 16'd24066;
          lut[1241] <= 16'd24085;
          lut[1242] <= 16'd24103;
          lut[1243] <= 16'd24121;
          lut[1244] <= 16'd24138;
          lut[1245] <= 16'd24155;
          lut[1246] <= 16'd24172;
          lut[1247] <= 16'd24188;
          lut[1248] <= 16'd24204;
          lut[1249] <= 16'd24220;
          lut[1250] <= 16'd24235;
          lut[1251] <= 16'd24251;
          lut[1252] <= 16'd24265;
          lut[1253] <= 16'd24280;
          lut[1254] <= 16'd24294;
          lut[1255] <= 16'd24308;
          lut[1256] <= 16'd24322;
          lut[1257] <= 16'd24335;
          lut[1258] <= 16'd24348;
          lut[1259] <= 16'd24361;
          lut[1260] <= 16'd24374;
          lut[1261] <= 16'd24386;
          lut[1262] <= 16'd24398;
          lut[1263] <= 16'd24410;
          lut[1264] <= 16'd24422;
          lut[1265] <= 16'd24434;
          lut[1266] <= 16'd24445;
          lut[1267] <= 16'd24456;
          lut[1268] <= 16'd24467;
          lut[1269] <= 16'd24478;
          lut[1270] <= 16'd24489;
          lut[1271] <= 16'd24499;
          lut[1272] <= 16'd24509;
          lut[1273] <= 16'd24520;
          lut[1274] <= 16'd24529;
          lut[1275] <= 16'd24539;
          lut[1276] <= 16'd24549;
          lut[1277] <= 16'd24558;
          lut[1278] <= 16'd24568;
          lut[1279] <= 16'd24577;
          lut[1280] <= 0;
          lut[1281] <= 16'd1633;
          lut[1282] <= 16'd3234;
          lut[1283] <= 16'd4775;
          lut[1284] <= 16'd6234;
          lut[1285] <= 16'd7596;
          lut[1286] <= 16'd8854;
          lut[1287] <= 16'd10006;
          lut[1288] <= 16'd11055;
          lut[1289] <= 16'd12006;
          lut[1290] <= 16'd12868;
          lut[1291] <= 16'd13648;
          lut[1292] <= 16'd14353;
          lut[1293] <= 16'd14993;
          lut[1294] <= 16'd15574;
          lut[1295] <= 16'd16102;
          lut[1296] <= 16'd16584;
          lut[1297] <= 16'd17024;
          lut[1298] <= 16'd17428;
          lut[1299] <= 16'd17798;
          lut[1300] <= 16'd18140;
          lut[1301] <= 16'd18455;
          lut[1302] <= 16'd18746;
          lut[1303] <= 16'd19016;
          lut[1304] <= 16'd19268;
          lut[1305] <= 16'd19502;
          lut[1306] <= 16'd19720;
          lut[1307] <= 16'd19924;
          lut[1308] <= 16'd20116;
          lut[1309] <= 16'd20295;
          lut[1310] <= 16'd20464;
          lut[1311] <= 16'd20623;
          lut[1312] <= 16'd20773;
          lut[1313] <= 16'd20915;
          lut[1314] <= 16'd21049;
          lut[1315] <= 16'd21176;
          lut[1316] <= 16'd21297;
          lut[1317] <= 16'd21411;
          lut[1318] <= 16'd21520;
          lut[1319] <= 16'd21623;
          lut[1320] <= 16'd21722;
          lut[1321] <= 16'd21816;
          lut[1322] <= 16'd21906;
          lut[1323] <= 16'd21992;
          lut[1324] <= 16'd22074;
          lut[1325] <= 16'd22153;
          lut[1326] <= 16'd22229;
          lut[1327] <= 16'd22301;
          lut[1328] <= 16'd22371;
          lut[1329] <= 16'd22438;
          lut[1330] <= 16'd22502;
          lut[1331] <= 16'd22564;
          lut[1332] <= 16'd22623;
          lut[1333] <= 16'd22681;
          lut[1334] <= 16'd22736;
          lut[1335] <= 16'd22789;
          lut[1336] <= 16'd22841;
          lut[1337] <= 16'd22890;
          lut[1338] <= 16'd22939;
          lut[1339] <= 16'd22985;
          lut[1340] <= 16'd23030;
          lut[1341] <= 16'd23074;
          lut[1342] <= 16'd23116;
          lut[1343] <= 16'd23157;
          lut[1344] <= 16'd23196;
          lut[1345] <= 16'd23235;
          lut[1346] <= 16'd23272;
          lut[1347] <= 16'd23308;
          lut[1348] <= 16'd23344;
          lut[1349] <= 16'd23378;
          lut[1350] <= 16'd23411;
          lut[1351] <= 16'd23443;
          lut[1352] <= 16'd23475;
          lut[1353] <= 16'd23505;
          lut[1354] <= 16'd23535;
          lut[1355] <= 16'd23564;
          lut[1356] <= 16'd23592;
          lut[1357] <= 16'd23620;
          lut[1358] <= 16'd23647;
          lut[1359] <= 16'd23673;
          lut[1360] <= 16'd23698;
          lut[1361] <= 16'd23723;
          lut[1362] <= 16'd23748;
          lut[1363] <= 16'd23771;
          lut[1364] <= 16'd23795;
          lut[1365] <= 16'd23817;
          lut[1366] <= 16'd23839;
          lut[1367] <= 16'd23861;
          lut[1368] <= 16'd23882;
          lut[1369] <= 16'd23903;
          lut[1370] <= 16'd23923;
          lut[1371] <= 16'd23943;
          lut[1372] <= 16'd23962;
          lut[1373] <= 16'd23981;
          lut[1374] <= 16'd23999;
          lut[1375] <= 16'd24018;
          lut[1376] <= 16'd24035;
          lut[1377] <= 16'd24053;
          lut[1378] <= 16'd24070;
          lut[1379] <= 16'd24087;
          lut[1380] <= 16'd24103;
          lut[1381] <= 16'd24119;
          lut[1382] <= 16'd24135;
          lut[1383] <= 16'd24150;
          lut[1384] <= 16'd24165;
          lut[1385] <= 16'd24180;
          lut[1386] <= 16'd24195;
          lut[1387] <= 16'd24209;
          lut[1388] <= 16'd24223;
          lut[1389] <= 16'd24237;
          lut[1390] <= 16'd24251;
          lut[1391] <= 16'd24264;
          lut[1392] <= 16'd24277;
          lut[1393] <= 16'd24290;
          lut[1394] <= 16'd24302;
          lut[1395] <= 16'd24315;
          lut[1396] <= 16'd24327;
          lut[1397] <= 16'd24339;
          lut[1398] <= 16'd24351;
          lut[1399] <= 16'd24362;
          lut[1400] <= 16'd24374;
          lut[1401] <= 16'd24385;
          lut[1402] <= 16'd24396;
          lut[1403] <= 16'd24407;
          lut[1404] <= 16'd24417;
          lut[1405] <= 16'd24428;
          lut[1406] <= 16'd24438;
          lut[1407] <= 16'd24449;
          lut[1408] <= 0;
          lut[1409] <= 16'd1485;
          lut[1410] <= 16'd2947;
          lut[1411] <= 16'd4362;
          lut[1412] <= 16'd5714;
          lut[1413] <= 16'd6990;
          lut[1414] <= 16'd8181;
          lut[1415] <= 16'd9285;
          lut[1416] <= 16'd10302;
          lut[1417] <= 16'd11235;
          lut[1418] <= 16'd12088;
          lut[1419] <= 16'd12868;
          lut[1420] <= 16'd13580;
          lut[1421] <= 16'd14230;
          lut[1422] <= 16'd14825;
          lut[1423] <= 16'd15369;
          lut[1424] <= 16'd15868;
          lut[1425] <= 16'd16327;
          lut[1426] <= 16'd16748;
          lut[1427] <= 16'd17138;
          lut[1428] <= 16'd17497;
          lut[1429] <= 16'd17830;
          lut[1430] <= 16'd18140;
          lut[1431] <= 16'd18427;
          lut[1432] <= 16'd18695;
          lut[1433] <= 16'd18945;
          lut[1434] <= 16'd19178;
          lut[1435] <= 16'd19397;
          lut[1436] <= 16'd19603;
          lut[1437] <= 16'd19796;
          lut[1438] <= 16'd19978;
          lut[1439] <= 16'd20149;
          lut[1440] <= 16'd20311;
          lut[1441] <= 16'd20464;
          lut[1442] <= 16'd20609;
          lut[1443] <= 16'd20747;
          lut[1444] <= 16'd20877;
          lut[1445] <= 16'd21001;
          lut[1446] <= 16'd21119;
          lut[1447] <= 16'd21232;
          lut[1448] <= 16'd21339;
          lut[1449] <= 16'd21441;
          lut[1450] <= 16'd21539;
          lut[1451] <= 16'd21633;
          lut[1452] <= 16'd21722;
          lut[1453] <= 16'd21808;
          lut[1454] <= 16'd21890;
          lut[1455] <= 16'd21969;
          lut[1456] <= 16'd22045;
          lut[1457] <= 16'd22118;
          lut[1458] <= 16'd22188;
          lut[1459] <= 16'd22255;
          lut[1460] <= 16'd22320;
          lut[1461] <= 16'd22383;
          lut[1462] <= 16'd22443;
          lut[1463] <= 16'd22502;
          lut[1464] <= 16'd22558;
          lut[1465] <= 16'd22612;
          lut[1466] <= 16'd22665;
          lut[1467] <= 16'd22716;
          lut[1468] <= 16'd22765;
          lut[1469] <= 16'd22813;
          lut[1470] <= 16'd22859;
          lut[1471] <= 16'd22904;
          lut[1472] <= 16'd22947;
          lut[1473] <= 16'd22989;
          lut[1474] <= 16'd23030;
          lut[1475] <= 16'd23070;
          lut[1476] <= 16'd23108;
          lut[1477] <= 16'd23146;
          lut[1478] <= 16'd23182;
          lut[1479] <= 16'd23218;
          lut[1480] <= 16'd23252;
          lut[1481] <= 16'd23286;
          lut[1482] <= 16'd23318;
          lut[1483] <= 16'd23350;
          lut[1484] <= 16'd23381;
          lut[1485] <= 16'd23411;
          lut[1486] <= 16'd23441;
          lut[1487] <= 16'd23469;
          lut[1488] <= 16'd23497;
          lut[1489] <= 16'd23524;
          lut[1490] <= 16'd23551;
          lut[1491] <= 16'd23577;
          lut[1492] <= 16'd23603;
          lut[1493] <= 16'd23627;
          lut[1494] <= 16'd23652;
          lut[1495] <= 16'd23675;
          lut[1496] <= 16'd23698;
          lut[1497] <= 16'd23721;
          lut[1498] <= 16'd23743;
          lut[1499] <= 16'd23765;
          lut[1500] <= 16'd23786;
          lut[1501] <= 16'd23807;
          lut[1502] <= 16'd23827;
          lut[1503] <= 16'd23847;
          lut[1504] <= 16'd23867;
          lut[1505] <= 16'd23886;
          lut[1506] <= 16'd23905;
          lut[1507] <= 16'd23923;
          lut[1508] <= 16'd23941;
          lut[1509] <= 16'd23959;
          lut[1510] <= 16'd23976;
          lut[1511] <= 16'd23993;
          lut[1512] <= 16'd24009;
          lut[1513] <= 16'd24026;
          lut[1514] <= 16'd24042;
          lut[1515] <= 16'd24057;
          lut[1516] <= 16'd24073;
          lut[1517] <= 16'd24088;
          lut[1518] <= 16'd24103;
          lut[1519] <= 16'd24118;
          lut[1520] <= 16'd24132;
          lut[1521] <= 16'd24146;
          lut[1522] <= 16'd24160;
          lut[1523] <= 16'd24174;
          lut[1524] <= 16'd24187;
          lut[1525] <= 16'd24200;
          lut[1526] <= 16'd24213;
          lut[1527] <= 16'd24226;
          lut[1528] <= 16'd24238;
          lut[1529] <= 16'd24251;
          lut[1530] <= 16'd24263;
          lut[1531] <= 16'd24275;
          lut[1532] <= 16'd24286;
          lut[1533] <= 16'd24298;
          lut[1534] <= 16'd24309;
          lut[1535] <= 16'd24320;
          lut[1536] <= 0;
          lut[1537] <= 16'd1362;
          lut[1538] <= 16'd2706;
          lut[1539] <= 16'd4014;
          lut[1540] <= 16'd5272;
          lut[1541] <= 16'd6468;
          lut[1542] <= 16'd7596;
          lut[1543] <= 16'd8652;
          lut[1544] <= 16'd9634;
          lut[1545] <= 16'd10543;
          lut[1546] <= 16'd11383;
          lut[1547] <= 16'd12156;
          lut[1548] <= 16'd12868;
          lut[1549] <= 16'd13523;
          lut[1550] <= 16'd14126;
          lut[1551] <= 16'd14681;
          lut[1552] <= 16'd15193;
          lut[1553] <= 16'd15665;
          lut[1554] <= 16'd16102;
          lut[1555] <= 16'd16507;
          lut[1556] <= 16'd16882;
          lut[1557] <= 16'd17230;
          lut[1558] <= 16'd17555;
          lut[1559] <= 16'd17857;
          lut[1560] <= 16'd18140;
          lut[1561] <= 16'd18404;
          lut[1562] <= 16'd18651;
          lut[1563] <= 16'd18884;
          lut[1564] <= 16'd19102;
          lut[1565] <= 16'd19308;
          lut[1566] <= 16'd19502;
          lut[1567] <= 16'd19685;
          lut[1568] <= 16'd19858;
          lut[1569] <= 16'd20022;
          lut[1570] <= 16'd20177;
          lut[1571] <= 16'd20324;
          lut[1572] <= 16'd20464;
          lut[1573] <= 16'd20598;
          lut[1574] <= 16'd20724;
          lut[1575] <= 16'd20845;
          lut[1576] <= 16'd20961;
          lut[1577] <= 16'd21071;
          lut[1578] <= 16'd21176;
          lut[1579] <= 16'd21277;
          lut[1580] <= 16'd21374;
          lut[1581] <= 16'd21466;
          lut[1582] <= 16'd21555;
          lut[1583] <= 16'd21640;
          lut[1584] <= 16'd21722;
          lut[1585] <= 16'd21801;
          lut[1586] <= 16'd21877;
          lut[1587] <= 16'd21950;
          lut[1588] <= 16'd22020;
          lut[1589] <= 16'd22088;
          lut[1590] <= 16'd22153;
          lut[1591] <= 16'd22216;
          lut[1592] <= 16'd22277;
          lut[1593] <= 16'd22336;
          lut[1594] <= 16'd22393;
          lut[1595] <= 16'd22448;
          lut[1596] <= 16'd22502;
          lut[1597] <= 16'd22553;
          lut[1598] <= 16'd22604;
          lut[1599] <= 16'd22652;
          lut[1600] <= 16'd22699;
          lut[1601] <= 16'd22745;
          lut[1602] <= 16'd22789;
          lut[1603] <= 16'd22832;
          lut[1604] <= 16'd22874;
          lut[1605] <= 16'd22915;
          lut[1606] <= 16'd22954;
          lut[1607] <= 16'd22993;
          lut[1608] <= 16'd23030;
          lut[1609] <= 16'd23067;
          lut[1610] <= 16'd23102;
          lut[1611] <= 16'd23137;
          lut[1612] <= 16'd23170;
          lut[1613] <= 16'd23203;
          lut[1614] <= 16'd23235;
          lut[1615] <= 16'd23266;
          lut[1616] <= 16'd23297;
          lut[1617] <= 16'd23326;
          lut[1618] <= 16'd23355;
          lut[1619] <= 16'd23383;
          lut[1620] <= 16'd23411;
          lut[1621] <= 16'd23438;
          lut[1622] <= 16'd23464;
          lut[1623] <= 16'd23490;
          lut[1624] <= 16'd23515;
          lut[1625] <= 16'd23540;
          lut[1626] <= 16'd23564;
          lut[1627] <= 16'd23588;
          lut[1628] <= 16'd23611;
          lut[1629] <= 16'd23633;
          lut[1630] <= 16'd23656;
          lut[1631] <= 16'd23677;
          lut[1632] <= 16'd23698;
          lut[1633] <= 16'd23719;
          lut[1634] <= 16'd23740;
          lut[1635] <= 16'd23760;
          lut[1636] <= 16'd23779;
          lut[1637] <= 16'd23798;
          lut[1638] <= 16'd23817;
          lut[1639] <= 16'd23836;
          lut[1640] <= 16'd23854;
          lut[1641] <= 16'd23872;
          lut[1642] <= 16'd23889;
          lut[1643] <= 16'd23906;
          lut[1644] <= 16'd23923;
          lut[1645] <= 16'd23939;
          lut[1646] <= 16'd23956;
          lut[1647] <= 16'd23972;
          lut[1648] <= 16'd23987;
          lut[1649] <= 16'd24003;
          lut[1650] <= 16'd24018;
          lut[1651] <= 16'd24032;
          lut[1652] <= 16'd24047;
          lut[1653] <= 16'd24061;
          lut[1654] <= 16'd24075;
          lut[1655] <= 16'd24089;
          lut[1656] <= 16'd24103;
          lut[1657] <= 16'd24116;
          lut[1658] <= 16'd24130;
          lut[1659] <= 16'd24143;
          lut[1660] <= 16'd24155;
          lut[1661] <= 16'd24168;
          lut[1662] <= 16'd24180;
          lut[1663] <= 16'd24192;
          lut[1664] <= 0;
          lut[1665] <= 16'd1258;
          lut[1666] <= 16'd2501;
          lut[1667] <= 16'd3716;
          lut[1668] <= 16'd4891;
          lut[1669] <= 16'd6016;
          lut[1670] <= 16'd7085;
          lut[1671] <= 16'd8093;
          lut[1672] <= 16'd9038;
          lut[1673] <= 16'd9921;
          lut[1674] <= 16'd10743;
          lut[1675] <= 16'd11506;
          lut[1676] <= 16'd12213;
          lut[1677] <= 16'd12868;
          lut[1678] <= 16'd13475;
          lut[1679] <= 16'd14036;
          lut[1680] <= 16'd14557;
          lut[1681] <= 16'd15040;
          lut[1682] <= 16'd15488;
          lut[1683] <= 16'd15905;
          lut[1684] <= 16'd16293;
          lut[1685] <= 16'd16654;
          lut[1686] <= 16'd16992;
          lut[1687] <= 16'd17307;
          lut[1688] <= 16'd17603;
          lut[1689] <= 16'd17879;
          lut[1690] <= 16'd18140;
          lut[1691] <= 16'd18384;
          lut[1692] <= 16'd18614;
          lut[1693] <= 16'd18831;
          lut[1694] <= 16'd19036;
          lut[1695] <= 16'd19230;
          lut[1696] <= 16'd19414;
          lut[1697] <= 16'd19587;
          lut[1698] <= 16'd19752;
          lut[1699] <= 16'd19909;
          lut[1700] <= 16'd20058;
          lut[1701] <= 16'd20200;
          lut[1702] <= 16'd20335;
          lut[1703] <= 16'd20464;
          lut[1704] <= 16'd20588;
          lut[1705] <= 16'd20705;
          lut[1706] <= 16'd20818;
          lut[1707] <= 16'd20926;
          lut[1708] <= 16'd21029;
          lut[1709] <= 16'd21128;
          lut[1710] <= 16'd21223;
          lut[1711] <= 16'd21315;
          lut[1712] <= 16'd21403;
          lut[1713] <= 16'd21487;
          lut[1714] <= 16'd21568;
          lut[1715] <= 16'd21647;
          lut[1716] <= 16'd21722;
          lut[1717] <= 16'd21795;
          lut[1718] <= 16'd21865;
          lut[1719] <= 16'd21933;
          lut[1720] <= 16'd21999;
          lut[1721] <= 16'd22062;
          lut[1722] <= 16'd22123;
          lut[1723] <= 16'd22183;
          lut[1724] <= 16'd22240;
          lut[1725] <= 16'd22296;
          lut[1726] <= 16'd22350;
          lut[1727] <= 16'd22402;
          lut[1728] <= 16'd22453;
          lut[1729] <= 16'd22502;
          lut[1730] <= 16'd22550;
          lut[1731] <= 16'd22596;
          lut[1732] <= 16'd22641;
          lut[1733] <= 16'd22685;
          lut[1734] <= 16'd22727;
          lut[1735] <= 16'd22769;
          lut[1736] <= 16'd22809;
          lut[1737] <= 16'd22848;
          lut[1738] <= 16'd22887;
          lut[1739] <= 16'd22924;
          lut[1740] <= 16'd22960;
          lut[1741] <= 16'd22996;
          lut[1742] <= 16'd23030;
          lut[1743] <= 16'd23064;
          lut[1744] <= 16'd23097;
          lut[1745] <= 16'd23129;
          lut[1746] <= 16'd23160;
          lut[1747] <= 16'd23190;
          lut[1748] <= 16'd23220;
          lut[1749] <= 16'd23249;
          lut[1750] <= 16'd23278;
          lut[1751] <= 16'd23306;
          lut[1752] <= 16'd23333;
          lut[1753] <= 16'd23360;
          lut[1754] <= 16'd23386;
          lut[1755] <= 16'd23411;
          lut[1756] <= 16'd23436;
          lut[1757] <= 16'd23460;
          lut[1758] <= 16'd23484;
          lut[1759] <= 16'd23508;
          lut[1760] <= 16'd23531;
          lut[1761] <= 16'd23553;
          lut[1762] <= 16'd23575;
          lut[1763] <= 16'd23597;
          lut[1764] <= 16'd23618;
          lut[1765] <= 16'd23639;
          lut[1766] <= 16'd23659;
          lut[1767] <= 16'd23679;
          lut[1768] <= 16'd23698;
          lut[1769] <= 16'd23718;
          lut[1770] <= 16'd23737;
          lut[1771] <= 16'd23755;
          lut[1772] <= 16'd23773;
          lut[1773] <= 16'd23791;
          lut[1774] <= 16'd23809;
          lut[1775] <= 16'd23826;
          lut[1776] <= 16'd23843;
          lut[1777] <= 16'd23859;
          lut[1778] <= 16'd23876;
          lut[1779] <= 16'd23892;
          lut[1780] <= 16'd23907;
          lut[1781] <= 16'd23923;
          lut[1782] <= 16'd23938;
          lut[1783] <= 16'd23953;
          lut[1784] <= 16'd23968;
          lut[1785] <= 16'd23982;
          lut[1786] <= 16'd23997;
          lut[1787] <= 16'd24011;
          lut[1788] <= 16'd24025;
          lut[1789] <= 16'd24038;
          lut[1790] <= 16'd24051;
          lut[1791] <= 16'd24065;
          lut[1792] <= 0;
          lut[1793] <= 16'd1168;
          lut[1794] <= 16'd2325;
          lut[1795] <= 16'd3459;
          lut[1796] <= 16'd4560;
          lut[1797] <= 16'd5620;
          lut[1798] <= 16'd6634;
          lut[1799] <= 16'd7596;
          lut[1800] <= 16'd8506;
          lut[1801] <= 16'd9361;
          lut[1802] <= 16'd10162;
          lut[1803] <= 16'd10911;
          lut[1804] <= 16'd11610;
          lut[1805] <= 16'd12261;
          lut[1806] <= 16'd12868;
          lut[1807] <= 16'd13433;
          lut[1808] <= 16'd13959;
          lut[1809] <= 16'd14449;
          lut[1810] <= 16'd14905;
          lut[1811] <= 16'd15332;
          lut[1812] <= 16'd15730;
          lut[1813] <= 16'd16102;
          lut[1814] <= 16'd16451;
          lut[1815] <= 16'd16777;
          lut[1816] <= 16'd17084;
          lut[1817] <= 16'd17372;
          lut[1818] <= 16'd17643;
          lut[1819] <= 16'd17899;
          lut[1820] <= 16'd18140;
          lut[1821] <= 16'd18367;
          lut[1822] <= 16'd18582;
          lut[1823] <= 16'd18786;
          lut[1824] <= 16'd18979;
          lut[1825] <= 16'd19162;
          lut[1826] <= 16'd19336;
          lut[1827] <= 16'd19502;
          lut[1828] <= 16'd19659;
          lut[1829] <= 16'd19809;
          lut[1830] <= 16'd19953;
          lut[1831] <= 16'd20089;
          lut[1832] <= 16'd20220;
          lut[1833] <= 16'd20345;
          lut[1834] <= 16'd20464;
          lut[1835] <= 16'd20579;
          lut[1836] <= 16'd20689;
          lut[1837] <= 16'd20794;
          lut[1838] <= 16'd20895;
          lut[1839] <= 16'd20993;
          lut[1840] <= 16'd21086;
          lut[1841] <= 16'd21176;
          lut[1842] <= 16'd21263;
          lut[1843] <= 16'd21346;
          lut[1844] <= 16'd21427;
          lut[1845] <= 16'd21505;
          lut[1846] <= 16'd21580;
          lut[1847] <= 16'd21652;
          lut[1848] <= 16'd21722;
          lut[1849] <= 16'd21790;
          lut[1850] <= 16'd21855;
          lut[1851] <= 16'd21919;
          lut[1852] <= 16'd21980;
          lut[1853] <= 16'd22040;
          lut[1854] <= 16'd22097;
          lut[1855] <= 16'd22153;
          lut[1856] <= 16'd22208;
          lut[1857] <= 16'd22260;
          lut[1858] <= 16'd22311;
          lut[1859] <= 16'd22361;
          lut[1860] <= 16'd22409;
          lut[1861] <= 16'd22456;
          lut[1862] <= 16'd22502;
          lut[1863] <= 16'd22546;
          lut[1864] <= 16'd22589;
          lut[1865] <= 16'd22631;
          lut[1866] <= 16'd22672;
          lut[1867] <= 16'd22712;
          lut[1868] <= 16'd22751;
          lut[1869] <= 16'd22789;
          lut[1870] <= 16'd22826;
          lut[1871] <= 16'd22862;
          lut[1872] <= 16'd22897;
          lut[1873] <= 16'd22932;
          lut[1874] <= 16'd22965;
          lut[1875] <= 16'd22998;
          lut[1876] <= 16'd23030;
          lut[1877] <= 16'd23061;
          lut[1878] <= 16'd23092;
          lut[1879] <= 16'd23122;
          lut[1880] <= 16'd23151;
          lut[1881] <= 16'd23180;
          lut[1882] <= 16'd23208;
          lut[1883] <= 16'd23235;
          lut[1884] <= 16'd23262;
          lut[1885] <= 16'd23288;
          lut[1886] <= 16'd23314;
          lut[1887] <= 16'd23339;
          lut[1888] <= 16'd23363;
          lut[1889] <= 16'd23387;
          lut[1890] <= 16'd23411;
          lut[1891] <= 16'd23434;
          lut[1892] <= 16'd23457;
          lut[1893] <= 16'd23479;
          lut[1894] <= 16'd23501;
          lut[1895] <= 16'd23523;
          lut[1896] <= 16'd23544;
          lut[1897] <= 16'd23564;
          lut[1898] <= 16'd23584;
          lut[1899] <= 16'd23604;
          lut[1900] <= 16'd23624;
          lut[1901] <= 16'd23643;
          lut[1902] <= 16'd23662;
          lut[1903] <= 16'd23680;
          lut[1904] <= 16'd23698;
          lut[1905] <= 16'd23716;
          lut[1906] <= 16'd23734;
          lut[1907] <= 16'd23751;
          lut[1908] <= 16'd23768;
          lut[1909] <= 16'd23785;
          lut[1910] <= 16'd23801;
          lut[1911] <= 16'd23817;
          lut[1912] <= 16'd23833;
          lut[1913] <= 16'd23849;
          lut[1914] <= 16'd23864;
          lut[1915] <= 16'd23879;
          lut[1916] <= 16'd23894;
          lut[1917] <= 16'd23909;
          lut[1918] <= 16'd23923;
          lut[1919] <= 16'd23937;
          lut[1920] <= 0;
          lut[1921] <= 16'd1091;
          lut[1922] <= 16'd2172;
          lut[1923] <= 16'd3234;
          lut[1924] <= 16'd4270;
          lut[1925] <= 16'd5272;
          lut[1926] <= 16'd6234;
          lut[1927] <= 16'd7154;
          lut[1928] <= 16'd8027;
          lut[1929] <= 16'd8854;
          lut[1930] <= 16'd9634;
          lut[1931] <= 16'd10367;
          lut[1932] <= 16'd11055;
          lut[1933] <= 16'd11700;
          lut[1934] <= 16'd12303;
          lut[1935] <= 16'd12868;
          lut[1936] <= 16'd13396;
          lut[1937] <= 16'd13891;
          lut[1938] <= 16'd14353;
          lut[1939] <= 16'd14787;
          lut[1940] <= 16'd15193;
          lut[1941] <= 16'd15574;
          lut[1942] <= 16'd15931;
          lut[1943] <= 16'd16268;
          lut[1944] <= 16'd16584;
          lut[1945] <= 16'd16882;
          lut[1946] <= 16'd17163;
          lut[1947] <= 16'd17428;
          lut[1948] <= 16'd17678;
          lut[1949] <= 16'd17915;
          lut[1950] <= 16'd18140;
          lut[1951] <= 16'd18352;
          lut[1952] <= 16'd18554;
          lut[1953] <= 16'd18746;
          lut[1954] <= 16'd18929;
          lut[1955] <= 16'd19102;
          lut[1956] <= 16'd19268;
          lut[1957] <= 16'd19426;
          lut[1958] <= 16'd19576;
          lut[1959] <= 16'd19720;
          lut[1960] <= 16'd19858;
          lut[1961] <= 16'd19990;
          lut[1962] <= 16'd20116;
          lut[1963] <= 16'd20237;
          lut[1964] <= 16'd20353;
          lut[1965] <= 16'd20464;
          lut[1966] <= 16'd20571;
          lut[1967] <= 16'd20674;
          lut[1968] <= 16'd20773;
          lut[1969] <= 16'd20869;
          lut[1970] <= 16'd20961;
          lut[1971] <= 16'd21049;
          lut[1972] <= 16'd21135;
          lut[1973] <= 16'd21217;
          lut[1974] <= 16'd21297;
          lut[1975] <= 16'd21374;
          lut[1976] <= 16'd21448;
          lut[1977] <= 16'd21520;
          lut[1978] <= 16'd21590;
          lut[1979] <= 16'd21657;
          lut[1980] <= 16'd21722;
          lut[1981] <= 16'd21785;
          lut[1982] <= 16'd21847;
          lut[1983] <= 16'd21906;
          lut[1984] <= 16'd21964;
          lut[1985] <= 16'd22020;
          lut[1986] <= 16'd22074;
          lut[1987] <= 16'd22127;
          lut[1988] <= 16'd22179;
          lut[1989] <= 16'd22229;
          lut[1990] <= 16'd22277;
          lut[1991] <= 16'd22325;
          lut[1992] <= 16'd22371;
          lut[1993] <= 16'd22416;
          lut[1994] <= 16'd22459;
          lut[1995] <= 16'd22502;
          lut[1996] <= 16'd22543;
          lut[1997] <= 16'd22584;
          lut[1998] <= 16'd22623;
          lut[1999] <= 16'd22662;
          lut[2000] <= 16'd22699;
          lut[2001] <= 16'd22736;
          lut[2002] <= 16'd22772;
          lut[2003] <= 16'd22807;
          lut[2004] <= 16'd22841;
          lut[2005] <= 16'd22874;
          lut[2006] <= 16'd22907;
          lut[2007] <= 16'd22939;
          lut[2008] <= 16'd22970;
          lut[2009] <= 16'd23000;
          lut[2010] <= 16'd23030;
          lut[2011] <= 16'd23059;
          lut[2012] <= 16'd23088;
          lut[2013] <= 16'd23116;
          lut[2014] <= 16'd23143;
          lut[2015] <= 16'd23170;
          lut[2016] <= 16'd23196;
          lut[2017] <= 16'd23222;
          lut[2018] <= 16'd23247;
          lut[2019] <= 16'd23272;
          lut[2020] <= 16'd23297;
          lut[2021] <= 16'd23320;
          lut[2022] <= 16'd23344;
          lut[2023] <= 16'd23367;
          lut[2024] <= 16'd23389;
          lut[2025] <= 16'd23411;
          lut[2026] <= 16'd23433;
          lut[2027] <= 16'd23454;
          lut[2028] <= 16'd23475;
          lut[2029] <= 16'd23495;
          lut[2030] <= 16'd23515;
          lut[2031] <= 16'd23535;
          lut[2032] <= 16'd23555;
          lut[2033] <= 16'd23574;
          lut[2034] <= 16'd23592;
          lut[2035] <= 16'd23611;
          lut[2036] <= 16'd23629;
          lut[2037] <= 16'd23647;
          lut[2038] <= 16'd23664;
          lut[2039] <= 16'd23682;
          lut[2040] <= 16'd23698;
          lut[2041] <= 16'd23715;
          lut[2042] <= 16'd23732;
          lut[2043] <= 16'd23748;
          lut[2044] <= 16'd23764;
          lut[2045] <= 16'd23779;
          lut[2046] <= 16'd23795;
          lut[2047] <= 16'd23810;
          lut[2048] <= 0;
          lut[2049] <= 16'd1023;
          lut[2050] <= 16'd2037;
          lut[2051] <= 16'd3037;
          lut[2052] <= 16'd4014;
          lut[2053] <= 16'd4962;
          lut[2054] <= 16'd5878;
          lut[2055] <= 16'd6757;
          lut[2056] <= 16'd7596;
          lut[2057] <= 16'd8395;
          lut[2058] <= 16'd9152;
          lut[2059] <= 16'd9868;
          lut[2060] <= 16'd10543;
          lut[2061] <= 16'd11179;
          lut[2062] <= 16'd11777;
          lut[2063] <= 16'd12340;
          lut[2064] <= 16'd12868;
          lut[2065] <= 16'd13364;
          lut[2066] <= 16'd13831;
          lut[2067] <= 16'd14269;
          lut[2068] <= 16'd14681;
          lut[2069] <= 16'd15069;
          lut[2070] <= 16'd15434;
          lut[2071] <= 16'd15778;
          lut[2072] <= 16'd16102;
          lut[2073] <= 16'd16408;
          lut[2074] <= 16'd16698;
          lut[2075] <= 16'd16971;
          lut[2076] <= 16'd17230;
          lut[2077] <= 16'd17476;
          lut[2078] <= 16'd17708;
          lut[2079] <= 16'd17929;
          lut[2080] <= 16'd18140;
          lut[2081] <= 16'd18339;
          lut[2082] <= 16'd18530;
          lut[2083] <= 16'd18711;
          lut[2084] <= 16'd18884;
          lut[2085] <= 16'd19049;
          lut[2086] <= 16'd19207;
          lut[2087] <= 16'd19357;
          lut[2088] <= 16'd19502;
          lut[2089] <= 16'd19640;
          lut[2090] <= 16'd19772;
          lut[2091] <= 16'd19900;
          lut[2092] <= 16'd20022;
          lut[2093] <= 16'd20139;
          lut[2094] <= 16'd20252;
          lut[2095] <= 16'd20360;
          lut[2096] <= 16'd20464;
          lut[2097] <= 16'd20565;
          lut[2098] <= 16'd20662;
          lut[2099] <= 16'd20755;
          lut[2100] <= 16'd20845;
          lut[2101] <= 16'd20932;
          lut[2102] <= 16'd21016;
          lut[2103] <= 16'd21098;
          lut[2104] <= 16'd21176;
          lut[2105] <= 16'd21252;
          lut[2106] <= 16'd21326;
          lut[2107] <= 16'd21397;
          lut[2108] <= 16'd21466;
          lut[2109] <= 16'd21533;
          lut[2110] <= 16'd21598;
          lut[2111] <= 16'd21661;
          lut[2112] <= 16'd21722;
          lut[2113] <= 16'd21782;
          lut[2114] <= 16'd21839;
          lut[2115] <= 16'd21895;
          lut[2116] <= 16'd21950;
          lut[2117] <= 16'd22003;
          lut[2118] <= 16'd22054;
          lut[2119] <= 16'd22104;
          lut[2120] <= 16'd22153;
          lut[2121] <= 16'd22201;
          lut[2122] <= 16'd22247;
          lut[2123] <= 16'd22292;
          lut[2124] <= 16'd22336;
          lut[2125] <= 16'd22379;
          lut[2126] <= 16'd22421;
          lut[2127] <= 16'd22462;
          lut[2128] <= 16'd22502;
          lut[2129] <= 16'd22541;
          lut[2130] <= 16'd22579;
          lut[2131] <= 16'd22616;
          lut[2132] <= 16'd22652;
          lut[2133] <= 16'd22688;
          lut[2134] <= 16'd22722;
          lut[2135] <= 16'd22756;
          lut[2136] <= 16'd22789;
          lut[2137] <= 16'd22822;
          lut[2138] <= 16'd22853;
          lut[2139] <= 16'd22884;
          lut[2140] <= 16'd22915;
          lut[2141] <= 16'd22945;
          lut[2142] <= 16'd22974;
          lut[2143] <= 16'd23002;
          lut[2144] <= 16'd23030;
          lut[2145] <= 16'd23058;
          lut[2146] <= 16'd23084;
          lut[2147] <= 16'd23111;
          lut[2148] <= 16'd23137;
          lut[2149] <= 16'd23162;
          lut[2150] <= 16'd23187;
          lut[2151] <= 16'd23211;
          lut[2152] <= 16'd23235;
          lut[2153] <= 16'd23258;
          lut[2154] <= 16'd23281;
          lut[2155] <= 16'd23304;
          lut[2156] <= 16'd23326;
          lut[2157] <= 16'd23348;
          lut[2158] <= 16'd23369;
          lut[2159] <= 16'd23390;
          lut[2160] <= 16'd23411;
          lut[2161] <= 16'd23431;
          lut[2162] <= 16'd23451;
          lut[2163] <= 16'd23471;
          lut[2164] <= 16'd23490;
          lut[2165] <= 16'd23509;
          lut[2166] <= 16'd23528;
          lut[2167] <= 16'd23546;
          lut[2168] <= 16'd23564;
          lut[2169] <= 16'd23582;
          lut[2170] <= 16'd23599;
          lut[2171] <= 16'd23617;
          lut[2172] <= 16'd23633;
          lut[2173] <= 16'd23650;
          lut[2174] <= 16'd23666;
          lut[2175] <= 16'd23683;
          lut[2176] <= 0;
          lut[2177] <= 16'd963;
          lut[2178] <= 16'd1919;
          lut[2179] <= 16'd2862;
          lut[2180] <= 16'd3786;
          lut[2181] <= 16'd4687;
          lut[2182] <= 16'd5559;
          lut[2183] <= 16'd6400;
          lut[2184] <= 16'd7206;
          lut[2185] <= 16'd7977;
          lut[2186] <= 16'd8712;
          lut[2187] <= 16'd9409;
          lut[2188] <= 16'd10071;
          lut[2189] <= 16'd10696;
          lut[2190] <= 16'd11287;
          lut[2191] <= 16'd11845;
          lut[2192] <= 16'd12372;
          lut[2193] <= 16'd12868;
          lut[2194] <= 16'd13336;
          lut[2195] <= 16'd13777;
          lut[2196] <= 16'd14193;
          lut[2197] <= 16'd14586;
          lut[2198] <= 16'd14957;
          lut[2199] <= 16'd15307;
          lut[2200] <= 16'd15639;
          lut[2201] <= 16'd15952;
          lut[2202] <= 16'd16248;
          lut[2203] <= 16'd16529;
          lut[2204] <= 16'd16796;
          lut[2205] <= 16'd17049;
          lut[2206] <= 16'd17289;
          lut[2207] <= 16'd17518;
          lut[2208] <= 16'd17735;
          lut[2209] <= 16'd17942;
          lut[2210] <= 16'd18140;
          lut[2211] <= 16'd18328;
          lut[2212] <= 16'd18508;
          lut[2213] <= 16'd18679;
          lut[2214] <= 16'd18844;
          lut[2215] <= 16'd19001;
          lut[2216] <= 16'd19152;
          lut[2217] <= 16'd19296;
          lut[2218] <= 16'd19435;
          lut[2219] <= 16'd19568;
          lut[2220] <= 16'd19695;
          lut[2221] <= 16'd19818;
          lut[2222] <= 16'd19936;
          lut[2223] <= 16'd20050;
          lut[2224] <= 16'd20159;
          lut[2225] <= 16'd20265;
          lut[2226] <= 16'd20366;
          lut[2227] <= 16'd20464;
          lut[2228] <= 16'd20559;
          lut[2229] <= 16'd20651;
          lut[2230] <= 16'd20739;
          lut[2231] <= 16'd20824;
          lut[2232] <= 16'd20907;
          lut[2233] <= 16'd20987;
          lut[2234] <= 16'd21065;
          lut[2235] <= 16'd21140;
          lut[2236] <= 16'd21212;
          lut[2237] <= 16'd21283;
          lut[2238] <= 16'd21351;
          lut[2239] <= 16'd21418;
          lut[2240] <= 16'd21482;
          lut[2241] <= 16'd21545;
          lut[2242] <= 16'd21606;
          lut[2243] <= 16'd21665;
          lut[2244] <= 16'd21722;
          lut[2245] <= 16'd21778;
          lut[2246] <= 16'd21833;
          lut[2247] <= 16'd21885;
          lut[2248] <= 16'd21937;
          lut[2249] <= 16'd21987;
          lut[2250] <= 16'd22036;
          lut[2251] <= 16'd22084;
          lut[2252] <= 16'd22130;
          lut[2253] <= 16'd22176;
          lut[2254] <= 16'd22220;
          lut[2255] <= 16'd22263;
          lut[2256] <= 16'd22305;
          lut[2257] <= 16'd22347;
          lut[2258] <= 16'd22387;
          lut[2259] <= 16'd22426;
          lut[2260] <= 16'd22464;
          lut[2261] <= 16'd22502;
          lut[2262] <= 16'd22538;
          lut[2263] <= 16'd22574;
          lut[2264] <= 16'd22609;
          lut[2265] <= 16'd22644;
          lut[2266] <= 16'd22677;
          lut[2267] <= 16'd22710;
          lut[2268] <= 16'd22742;
          lut[2269] <= 16'd22774;
          lut[2270] <= 16'd22805;
          lut[2271] <= 16'd22835;
          lut[2272] <= 16'd22864;
          lut[2273] <= 16'd22893;
          lut[2274] <= 16'd22922;
          lut[2275] <= 16'd22950;
          lut[2276] <= 16'd22977;
          lut[2277] <= 16'd23004;
          lut[2278] <= 16'd23030;
          lut[2279] <= 16'd23056;
          lut[2280] <= 16'd23081;
          lut[2281] <= 16'd23106;
          lut[2282] <= 16'd23130;
          lut[2283] <= 16'd23154;
          lut[2284] <= 16'd23178;
          lut[2285] <= 16'd23201;
          lut[2286] <= 16'd23224;
          lut[2287] <= 16'd23246;
          lut[2288] <= 16'd23268;
          lut[2289] <= 16'd23289;
          lut[2290] <= 16'd23311;
          lut[2291] <= 16'd23331;
          lut[2292] <= 16'd23352;
          lut[2293] <= 16'd23372;
          lut[2294] <= 16'd23392;
          lut[2295] <= 16'd23411;
          lut[2296] <= 16'd23430;
          lut[2297] <= 16'd23449;
          lut[2298] <= 16'd23468;
          lut[2299] <= 16'd23486;
          lut[2300] <= 16'd23504;
          lut[2301] <= 16'd23521;
          lut[2302] <= 16'd23539;
          lut[2303] <= 16'd23556;
          lut[2304] <= 0;
          lut[2305] <= 16'd909;
          lut[2306] <= 16'd1813;
          lut[2307] <= 16'd2706;
          lut[2308] <= 16'd3583;
          lut[2309] <= 16'd4439;
          lut[2310] <= 16'd5272;
          lut[2311] <= 16'd6077;
          lut[2312] <= 16'd6852;
          lut[2313] <= 16'd7596;
          lut[2314] <= 16'd8308;
          lut[2315] <= 16'd8987;
          lut[2316] <= 16'd9634;
          lut[2317] <= 16'd10248;
          lut[2318] <= 16'd10831;
          lut[2319] <= 16'd11383;
          lut[2320] <= 16'd11905;
          lut[2321] <= 16'd12400;
          lut[2322] <= 16'd12868;
          lut[2323] <= 16'd13311;
          lut[2324] <= 16'd13729;
          lut[2325] <= 16'd14126;
          lut[2326] <= 16'd14501;
          lut[2327] <= 16'd14856;
          lut[2328] <= 16'd15193;
          lut[2329] <= 16'd15512;
          lut[2330] <= 16'd15815;
          lut[2331] <= 16'd16102;
          lut[2332] <= 16'd16375;
          lut[2333] <= 16'd16635;
          lut[2334] <= 16'd16882;
          lut[2335] <= 16'd17117;
          lut[2336] <= 16'd17341;
          lut[2337] <= 16'd17555;
          lut[2338] <= 16'd17759;
          lut[2339] <= 16'd17953;
          lut[2340] <= 16'd18140;
          lut[2341] <= 16'd18318;
          lut[2342] <= 16'd18488;
          lut[2343] <= 16'd18651;
          lut[2344] <= 16'd18808;
          lut[2345] <= 16'd18958;
          lut[2346] <= 16'd19102;
          lut[2347] <= 16'd19241;
          lut[2348] <= 16'd19374;
          lut[2349] <= 16'd19502;
          lut[2350] <= 16'd19625;
          lut[2351] <= 16'd19744;
          lut[2352] <= 16'd19858;
          lut[2353] <= 16'd19968;
          lut[2354] <= 16'd20074;
          lut[2355] <= 16'd20177;
          lut[2356] <= 16'd20276;
          lut[2357] <= 16'd20372;
          lut[2358] <= 16'd20464;
          lut[2359] <= 16'd20554;
          lut[2360] <= 16'd20641;
          lut[2361] <= 16'd20724;
          lut[2362] <= 16'd20806;
          lut[2363] <= 16'd20884;
          lut[2364] <= 16'd20961;
          lut[2365] <= 16'd21035;
          lut[2366] <= 16'd21107;
          lut[2367] <= 16'd21176;
          lut[2368] <= 16'd21244;
          lut[2369] <= 16'd21310;
          lut[2370] <= 16'd21374;
          lut[2371] <= 16'd21436;
          lut[2372] <= 16'd21496;
          lut[2373] <= 16'd21555;
          lut[2374] <= 16'd21612;
          lut[2375] <= 16'd21668;
          lut[2376] <= 16'd21722;
          lut[2377] <= 16'd21775;
          lut[2378] <= 16'd21827;
          lut[2379] <= 16'd21877;
          lut[2380] <= 16'd21926;
          lut[2381] <= 16'd21973;
          lut[2382] <= 16'd22020;
          lut[2383] <= 16'd22066;
          lut[2384] <= 16'd22110;
          lut[2385] <= 16'd22153;
          lut[2386] <= 16'd22196;
          lut[2387] <= 16'd22237;
          lut[2388] <= 16'd22277;
          lut[2389] <= 16'd22317;
          lut[2390] <= 16'd22356;
          lut[2391] <= 16'd22393;
          lut[2392] <= 16'd22430;
          lut[2393] <= 16'd22466;
          lut[2394] <= 16'd22502;
          lut[2395] <= 16'd22536;
          lut[2396] <= 16'd22570;
          lut[2397] <= 16'd22604;
          lut[2398] <= 16'd22636;
          lut[2399] <= 16'd22668;
          lut[2400] <= 16'd22699;
          lut[2401] <= 16'd22730;
          lut[2402] <= 16'd22760;
          lut[2403] <= 16'd22789;
          lut[2404] <= 16'd22818;
          lut[2405] <= 16'd22846;
          lut[2406] <= 16'd22874;
          lut[2407] <= 16'd22901;
          lut[2408] <= 16'd22928;
          lut[2409] <= 16'd22954;
          lut[2410] <= 16'd22980;
          lut[2411] <= 16'd23005;
          lut[2412] <= 16'd23030;
          lut[2413] <= 16'd23055;
          lut[2414] <= 16'd23078;
          lut[2415] <= 16'd23102;
          lut[2416] <= 16'd23125;
          lut[2417] <= 16'd23148;
          lut[2418] <= 16'd23170;
          lut[2419] <= 16'd23192;
          lut[2420] <= 16'd23214;
          lut[2421] <= 16'd23235;
          lut[2422] <= 16'd23256;
          lut[2423] <= 16'd23276;
          lut[2424] <= 16'd23297;
          lut[2425] <= 16'd23316;
          lut[2426] <= 16'd23336;
          lut[2427] <= 16'd23355;
          lut[2428] <= 16'd23374;
          lut[2429] <= 16'd23393;
          lut[2430] <= 16'd23411;
          lut[2431] <= 16'd23429;
          lut[2432] <= 0;
          lut[2433] <= 16'd862;
          lut[2434] <= 16'd1718;
          lut[2435] <= 16'd2566;
          lut[2436] <= 16'd3400;
          lut[2437] <= 16'd4216;
          lut[2438] <= 16'd5012;
          lut[2439] <= 16'd5783;
          lut[2440] <= 16'd6529;
          lut[2441] <= 16'd7248;
          lut[2442] <= 16'd7938;
          lut[2443] <= 16'd8598;
          lut[2444] <= 16'd9229;
          lut[2445] <= 16'd9831;
          lut[2446] <= 16'd10404;
          lut[2447] <= 16'd10949;
          lut[2448] <= 16'd11467;
          lut[2449] <= 16'd11959;
          lut[2450] <= 16'd12425;
          lut[2451] <= 16'd12868;
          lut[2452] <= 16'd13288;
          lut[2453] <= 16'd13686;
          lut[2454] <= 16'd14065;
          lut[2455] <= 16'd14424;
          lut[2456] <= 16'd14765;
          lut[2457] <= 16'd15088;
          lut[2458] <= 16'd15396;
          lut[2459] <= 16'd15689;
          lut[2460] <= 16'd15968;
          lut[2461] <= 16'd16233;
          lut[2462] <= 16'd16486;
          lut[2463] <= 16'd16727;
          lut[2464] <= 16'd16957;
          lut[2465] <= 16'd17177;
          lut[2466] <= 16'd17387;
          lut[2467] <= 16'd17587;
          lut[2468] <= 16'd17779;
          lut[2469] <= 16'd17963;
          lut[2470] <= 16'd18140;
          lut[2471] <= 16'd18308;
          lut[2472] <= 16'd18470;
          lut[2473] <= 16'd18626;
          lut[2474] <= 16'd18775;
          lut[2475] <= 16'd18919;
          lut[2476] <= 16'd19057;
          lut[2477] <= 16'd19190;
          lut[2478] <= 16'd19318;
          lut[2479] <= 16'd19442;
          lut[2480] <= 16'd19561;
          lut[2481] <= 16'd19675;
          lut[2482] <= 16'd19786;
          lut[2483] <= 16'd19893;
          lut[2484] <= 16'd19996;
          lut[2485] <= 16'd20096;
          lut[2486] <= 16'd20193;
          lut[2487] <= 16'd20286;
          lut[2488] <= 16'd20377;
          lut[2489] <= 16'd20464;
          lut[2490] <= 16'd20549;
          lut[2491] <= 16'd20632;
          lut[2492] <= 16'd20711;
          lut[2493] <= 16'd20789;
          lut[2494] <= 16'd20864;
          lut[2495] <= 16'd20937;
          lut[2496] <= 16'd21008;
          lut[2497] <= 16'd21077;
          lut[2498] <= 16'd21143;
          lut[2499] <= 16'd21209;
          lut[2500] <= 16'd21272;
          lut[2501] <= 16'd21333;
          lut[2502] <= 16'd21393;
          lut[2503] <= 16'd21452;
          lut[2504] <= 16'd21509;
          lut[2505] <= 16'd21564;
          lut[2506] <= 16'd21618;
          lut[2507] <= 16'd21671;
          lut[2508] <= 16'd21722;
          lut[2509] <= 16'd21772;
          lut[2510] <= 16'd21821;
          lut[2511] <= 16'd21869;
          lut[2512] <= 16'd21916;
          lut[2513] <= 16'd21961;
          lut[2514] <= 16'd22005;
          lut[2515] <= 16'd22049;
          lut[2516] <= 16'd22091;
          lut[2517] <= 16'd22133;
          lut[2518] <= 16'd22173;
          lut[2519] <= 16'd22213;
          lut[2520] <= 16'd22252;
          lut[2521] <= 16'd22290;
          lut[2522] <= 16'd22327;
          lut[2523] <= 16'd22364;
          lut[2524] <= 16'd22399;
          lut[2525] <= 16'd22434;
          lut[2526] <= 16'd22468;
          lut[2527] <= 16'd22502;
          lut[2528] <= 16'd22535;
          lut[2529] <= 16'd22567;
          lut[2530] <= 16'd22598;
          lut[2531] <= 16'd22629;
          lut[2532] <= 16'd22660;
          lut[2533] <= 16'd22689;
          lut[2534] <= 16'd22719;
          lut[2535] <= 16'd22747;
          lut[2536] <= 16'd22775;
          lut[2537] <= 16'd22803;
          lut[2538] <= 16'd22830;
          lut[2539] <= 16'd22857;
          lut[2540] <= 16'd22883;
          lut[2541] <= 16'd22908;
          lut[2542] <= 16'd22934;
          lut[2543] <= 16'd22958;
          lut[2544] <= 16'd22983;
          lut[2545] <= 16'd23007;
          lut[2546] <= 16'd23030;
          lut[2547] <= 16'd23053;
          lut[2548] <= 16'd23076;
          lut[2549] <= 16'd23098;
          lut[2550] <= 16'd23120;
          lut[2551] <= 16'd23142;
          lut[2552] <= 16'd23163;
          lut[2553] <= 16'd23184;
          lut[2554] <= 16'd23205;
          lut[2555] <= 16'd23225;
          lut[2556] <= 16'd23245;
          lut[2557] <= 16'd23264;
          lut[2558] <= 16'd23284;
          lut[2559] <= 16'd23303;
          lut[2560] <= 0;
          lut[2561] <= 16'd819;
          lut[2562] <= 16'd1633;
          lut[2563] <= 16'd2439;
          lut[2564] <= 16'd3234;
          lut[2565] <= 16'd4014;
          lut[2566] <= 16'd4775;
          lut[2567] <= 16'd5516;
          lut[2568] <= 16'd6234;
          lut[2569] <= 16'd6928;
          lut[2570] <= 16'd7596;
          lut[2571] <= 16'd8239;
          lut[2572] <= 16'd8854;
          lut[2573] <= 16'd9443;
          lut[2574] <= 16'd10006;
          lut[2575] <= 16'd10543;
          lut[2576] <= 16'd11055;
          lut[2577] <= 16'd11542;
          lut[2578] <= 16'd12006;
          lut[2579] <= 16'd12448;
          lut[2580] <= 16'd12868;
          lut[2581] <= 16'd13267;
          lut[2582] <= 16'd13648;
          lut[2583] <= 16'd14009;
          lut[2584] <= 16'd14353;
          lut[2585] <= 16'd14681;
          lut[2586] <= 16'd14993;
          lut[2587] <= 16'd15290;
          lut[2588] <= 16'd15574;
          lut[2589] <= 16'd15844;
          lut[2590] <= 16'd16102;
          lut[2591] <= 16'd16348;
          lut[2592] <= 16'd16584;
          lut[2593] <= 16'd16809;
          lut[2594] <= 16'd17024;
          lut[2595] <= 16'd17230;
          lut[2596] <= 16'd17428;
          lut[2597] <= 16'd17617;
          lut[2598] <= 16'd17798;
          lut[2599] <= 16'd17972;
          lut[2600] <= 16'd18140;
          lut[2601] <= 16'd18300;
          lut[2602] <= 16'd18455;
          lut[2603] <= 16'd18603;
          lut[2604] <= 16'd18746;
          lut[2605] <= 16'd18884;
          lut[2606] <= 16'd19016;
          lut[2607] <= 16'd19144;
          lut[2608] <= 16'd19268;
          lut[2609] <= 16'd19387;
          lut[2610] <= 16'd19502;
          lut[2611] <= 16'd19613;
          lut[2612] <= 16'd19720;
          lut[2613] <= 16'd19824;
          lut[2614] <= 16'd19924;
          lut[2615] <= 16'd20022;
          lut[2616] <= 16'd20116;
          lut[2617] <= 16'd20207;
          lut[2618] <= 16'd20295;
          lut[2619] <= 16'd20381;
          lut[2620] <= 16'd20464;
          lut[2621] <= 16'd20545;
          lut[2622] <= 16'd20623;
          lut[2623] <= 16'd20700;
          lut[2624] <= 16'd20773;
          lut[2625] <= 16'd20845;
          lut[2626] <= 16'd20915;
          lut[2627] <= 16'd20983;
          lut[2628] <= 16'd21049;
          lut[2629] <= 16'd21114;
          lut[2630] <= 16'd21176;
          lut[2631] <= 16'd21237;
          lut[2632] <= 16'd21297;
          lut[2633] <= 16'd21355;
          lut[2634] <= 16'd21411;
          lut[2635] <= 16'd21466;
          lut[2636] <= 16'd21520;
          lut[2637] <= 16'd21572;
          lut[2638] <= 16'd21623;
          lut[2639] <= 16'd21673;
          lut[2640] <= 16'd21722;
          lut[2641] <= 16'd21770;
          lut[2642] <= 16'd21816;
          lut[2643] <= 16'd21862;
          lut[2644] <= 16'd21906;
          lut[2645] <= 16'd21950;
          lut[2646] <= 16'd21992;
          lut[2647] <= 16'd22034;
          lut[2648] <= 16'd22074;
          lut[2649] <= 16'd22114;
          lut[2650] <= 16'd22153;
          lut[2651] <= 16'd22191;
          lut[2652] <= 16'd22229;
          lut[2653] <= 16'd22265;
          lut[2654] <= 16'd22301;
          lut[2655] <= 16'd22336;
          lut[2656] <= 16'd22371;
          lut[2657] <= 16'd22404;
          lut[2658] <= 16'd22438;
          lut[2659] <= 16'd22470;
          lut[2660] <= 16'd22502;
          lut[2661] <= 16'd22533;
          lut[2662] <= 16'd22564;
          lut[2663] <= 16'd22594;
          lut[2664] <= 16'd22623;
          lut[2665] <= 16'd22652;
          lut[2666] <= 16'd22681;
          lut[2667] <= 16'd22708;
          lut[2668] <= 16'd22736;
          lut[2669] <= 16'd22763;
          lut[2670] <= 16'd22789;
          lut[2671] <= 16'd22815;
          lut[2672] <= 16'd22841;
          lut[2673] <= 16'd22866;
          lut[2674] <= 16'd22890;
          lut[2675] <= 16'd22915;
          lut[2676] <= 16'd22939;
          lut[2677] <= 16'd22962;
          lut[2678] <= 16'd22985;
          lut[2679] <= 16'd23008;
          lut[2680] <= 16'd23030;
          lut[2681] <= 16'd23052;
          lut[2682] <= 16'd23074;
          lut[2683] <= 16'd23095;
          lut[2684] <= 16'd23116;
          lut[2685] <= 16'd23137;
          lut[2686] <= 16'd23157;
          lut[2687] <= 16'd23177;
          lut[2688] <= 0;
          lut[2689] <= 16'd780;
          lut[2690] <= 16'd1556;
          lut[2691] <= 16'd2325;
          lut[2692] <= 16'd3084;
          lut[2693] <= 16'd3830;
          lut[2694] <= 16'd4560;
          lut[2695] <= 16'd5272;
          lut[2696] <= 16'd5963;
          lut[2697] <= 16'd6634;
          lut[2698] <= 16'd7281;
          lut[2699] <= 16'd7905;
          lut[2700] <= 16'd8506;
          lut[2701] <= 16'd9082;
          lut[2702] <= 16'd9634;
          lut[2703] <= 16'd10162;
          lut[2704] <= 16'd10667;
          lut[2705] <= 16'd11150;
          lut[2706] <= 16'd11610;
          lut[2707] <= 16'd12049;
          lut[2708] <= 16'd12468;
          lut[2709] <= 16'd12868;
          lut[2710] <= 16'd13249;
          lut[2711] <= 16'd13612;
          lut[2712] <= 16'd13959;
          lut[2713] <= 16'd14289;
          lut[2714] <= 16'd14604;
          lut[2715] <= 16'd14905;
          lut[2716] <= 16'd15193;
          lut[2717] <= 16'd15467;
          lut[2718] <= 16'd15730;
          lut[2719] <= 16'd15981;
          lut[2720] <= 16'd16221;
          lut[2721] <= 16'd16451;
          lut[2722] <= 16'd16671;
          lut[2723] <= 16'd16882;
          lut[2724] <= 16'd17084;
          lut[2725] <= 16'd17278;
          lut[2726] <= 16'd17464;
          lut[2727] <= 16'd17643;
          lut[2728] <= 16'd17815;
          lut[2729] <= 16'd17980;
          lut[2730] <= 16'd18140;
          lut[2731] <= 16'd18293;
          lut[2732] <= 16'd18440;
          lut[2733] <= 16'd18582;
          lut[2734] <= 16'd18719;
          lut[2735] <= 16'd18851;
          lut[2736] <= 16'd18979;
          lut[2737] <= 16'd19102;
          lut[2738] <= 16'd19221;
          lut[2739] <= 16'd19336;
          lut[2740] <= 16'd19447;
          lut[2741] <= 16'd19555;
          lut[2742] <= 16'd19659;
          lut[2743] <= 16'd19760;
          lut[2744] <= 16'd19858;
          lut[2745] <= 16'd19953;
          lut[2746] <= 16'd20044;
          lut[2747] <= 16'd20133;
          lut[2748] <= 16'd20220;
          lut[2749] <= 16'd20304;
          lut[2750] <= 16'd20385;
          lut[2751] <= 16'd20464;
          lut[2752] <= 16'd20541;
          lut[2753] <= 16'd20616;
          lut[2754] <= 16'd20689;
          lut[2755] <= 16'd20760;
          lut[2756] <= 16'd20828;
          lut[2757] <= 16'd20895;
          lut[2758] <= 16'd20961;
          lut[2759] <= 16'd21024;
          lut[2760] <= 16'd21086;
          lut[2761] <= 16'd21147;
          lut[2762] <= 16'd21206;
          lut[2763] <= 16'd21263;
          lut[2764] <= 16'd21319;
          lut[2765] <= 16'd21374;
          lut[2766] <= 16'd21427;
          lut[2767] <= 16'd21479;
          lut[2768] <= 16'd21530;
          lut[2769] <= 16'd21580;
          lut[2770] <= 16'd21628;
          lut[2771] <= 16'd21676;
          lut[2772] <= 16'd21722;
          lut[2773] <= 16'd21768;
          lut[2774] <= 16'd21812;
          lut[2775] <= 16'd21855;
          lut[2776] <= 16'd21898;
          lut[2777] <= 16'd21939;
          lut[2778] <= 16'd21980;
          lut[2779] <= 16'd22020;
          lut[2780] <= 16'd22059;
          lut[2781] <= 16'd22097;
          lut[2782] <= 16'd22135;
          lut[2783] <= 16'd22172;
          lut[2784] <= 16'd22208;
          lut[2785] <= 16'd22243;
          lut[2786] <= 16'd22277;
          lut[2787] <= 16'd22311;
          lut[2788] <= 16'd22345;
          lut[2789] <= 16'd22377;
          lut[2790] <= 16'd22409;
          lut[2791] <= 16'd22441;
          lut[2792] <= 16'd22472;
          lut[2793] <= 16'd22502;
          lut[2794] <= 16'd22532;
          lut[2795] <= 16'd22561;
          lut[2796] <= 16'd22589;
          lut[2797] <= 16'd22618;
          lut[2798] <= 16'd22645;
          lut[2799] <= 16'd22672;
          lut[2800] <= 16'd22699;
          lut[2801] <= 16'd22725;
          lut[2802] <= 16'd22751;
          lut[2803] <= 16'd22777;
          lut[2804] <= 16'd22802;
          lut[2805] <= 16'd22826;
          lut[2806] <= 16'd22850;
          lut[2807] <= 16'd22874;
          lut[2808] <= 16'd22897;
          lut[2809] <= 16'd22920;
          lut[2810] <= 16'd22943;
          lut[2811] <= 16'd22965;
          lut[2812] <= 16'd22987;
          lut[2813] <= 16'd23009;
          lut[2814] <= 16'd23030;
          lut[2815] <= 16'd23051;
          lut[2816] <= 0;
          lut[2817] <= 16'd744;
          lut[2818] <= 16'd1485;
          lut[2819] <= 16'd2220;
          lut[2820] <= 16'd2947;
          lut[2821] <= 16'd3661;
          lut[2822] <= 16'd4362;
          lut[2823] <= 16'd5047;
          lut[2824] <= 16'd5714;
          lut[2825] <= 16'd6362;
          lut[2826] <= 16'd6990;
          lut[2827] <= 16'd7596;
          lut[2828] <= 16'd8181;
          lut[2829] <= 16'd8744;
          lut[2830] <= 16'd9285;
          lut[2831] <= 16'd9804;
          lut[2832] <= 16'd10302;
          lut[2833] <= 16'd10779;
          lut[2834] <= 16'd11235;
          lut[2835] <= 16'd11671;
          lut[2836] <= 16'd12088;
          lut[2837] <= 16'd12487;
          lut[2838] <= 16'd12868;
          lut[2839] <= 16'd13232;
          lut[2840] <= 16'd13580;
          lut[2841] <= 16'd13912;
          lut[2842] <= 16'd14230;
          lut[2843] <= 16'd14534;
          lut[2844] <= 16'd14825;
          lut[2845] <= 16'd15103;
          lut[2846] <= 16'd15369;
          lut[2847] <= 16'd15624;
          lut[2848] <= 16'd15868;
          lut[2849] <= 16'd16102;
          lut[2850] <= 16'd16327;
          lut[2851] <= 16'd16542;
          lut[2852] <= 16'd16748;
          lut[2853] <= 16'd16947;
          lut[2854] <= 16'd17138;
          lut[2855] <= 16'd17321;
          lut[2856] <= 16'd17497;
          lut[2857] <= 16'd17667;
          lut[2858] <= 16'd17830;
          lut[2859] <= 16'd17988;
          lut[2860] <= 16'd18140;
          lut[2861] <= 16'd18286;
          lut[2862] <= 16'd18427;
          lut[2863] <= 16'd18563;
          lut[2864] <= 16'd18695;
          lut[2865] <= 16'd18822;
          lut[2866] <= 16'd18945;
          lut[2867] <= 16'd19063;
          lut[2868] <= 16'd19178;
          lut[2869] <= 16'd19290;
          lut[2870] <= 16'd19397;
          lut[2871] <= 16'd19502;
          lut[2872] <= 16'd19603;
          lut[2873] <= 16'd19701;
          lut[2874] <= 16'd19796;
          lut[2875] <= 16'd19888;
          lut[2876] <= 16'd19978;
          lut[2877] <= 16'd20065;
          lut[2878] <= 16'd20149;
          lut[2879] <= 16'd20231;
          lut[2880] <= 16'd20311;
          lut[2881] <= 16'd20389;
          lut[2882] <= 16'd20464;
          lut[2883] <= 16'd20538;
          lut[2884] <= 16'd20609;
          lut[2885] <= 16'd20679;
          lut[2886] <= 16'd20747;
          lut[2887] <= 16'd20813;
          lut[2888] <= 16'd20877;
          lut[2889] <= 16'd20940;
          lut[2890] <= 16'd21001;
          lut[2891] <= 16'd21061;
          lut[2892] <= 16'd21119;
          lut[2893] <= 16'd21176;
          lut[2894] <= 16'd21232;
          lut[2895] <= 16'd21286;
          lut[2896] <= 16'd21339;
          lut[2897] <= 16'd21391;
          lut[2898] <= 16'd21441;
          lut[2899] <= 16'd21491;
          lut[2900] <= 16'd21539;
          lut[2901] <= 16'd21586;
          lut[2902] <= 16'd21633;
          lut[2903] <= 16'd21678;
          lut[2904] <= 16'd21722;
          lut[2905] <= 16'd21766;
          lut[2906] <= 16'd21808;
          lut[2907] <= 16'd21850;
          lut[2908] <= 16'd21890;
          lut[2909] <= 16'd21930;
          lut[2910] <= 16'd21969;
          lut[2911] <= 16'd22007;
          lut[2912] <= 16'd22045;
          lut[2913] <= 16'd22082;
          lut[2914] <= 16'd22118;
          lut[2915] <= 16'd22153;
          lut[2916] <= 16'd22188;
          lut[2917] <= 16'd22222;
          lut[2918] <= 16'd22255;
          lut[2919] <= 16'd22288;
          lut[2920] <= 16'd22320;
          lut[2921] <= 16'd22352;
          lut[2922] <= 16'd22383;
          lut[2923] <= 16'd22414;
          lut[2924] <= 16'd22443;
          lut[2925] <= 16'd22473;
          lut[2926] <= 16'd22502;
          lut[2927] <= 16'd22530;
          lut[2928] <= 16'd22558;
          lut[2929] <= 16'd22586;
          lut[2930] <= 16'd22612;
          lut[2931] <= 16'd22639;
          lut[2932] <= 16'd22665;
          lut[2933] <= 16'd22691;
          lut[2934] <= 16'd22716;
          lut[2935] <= 16'd22741;
          lut[2936] <= 16'd22765;
          lut[2937] <= 16'd22789;
          lut[2938] <= 16'd22813;
          lut[2939] <= 16'd22836;
          lut[2940] <= 16'd22859;
          lut[2941] <= 16'd22882;
          lut[2942] <= 16'd22904;
          lut[2943] <= 16'd22926;
          lut[2944] <= 0;
          lut[2945] <= 16'd712;
          lut[2946] <= 16'd1421;
          lut[2947] <= 16'd2125;
          lut[2948] <= 16'd2821;
          lut[2949] <= 16'd3507;
          lut[2950] <= 16'd4181;
          lut[2951] <= 16'd4841;
          lut[2952] <= 16'd5484;
          lut[2953] <= 16'd6111;
          lut[2954] <= 16'd6720;
          lut[2955] <= 16'd7309;
          lut[2956] <= 16'd7879;
          lut[2957] <= 16'd8429;
          lut[2958] <= 16'd8959;
          lut[2959] <= 16'd9468;
          lut[2960] <= 16'd9958;
          lut[2961] <= 16'd10429;
          lut[2962] <= 16'd10880;
          lut[2963] <= 16'd11312;
          lut[2964] <= 16'd11727;
          lut[2965] <= 16'd12124;
          lut[2966] <= 16'd12504;
          lut[2967] <= 16'd12868;
          lut[2968] <= 16'd13217;
          lut[2969] <= 16'd13550;
          lut[2970] <= 16'd13870;
          lut[2971] <= 16'd14176;
          lut[2972] <= 16'd14469;
          lut[2973] <= 16'd14750;
          lut[2974] <= 16'd15019;
          lut[2975] <= 16'd15278;
          lut[2976] <= 16'd15525;
          lut[2977] <= 16'd15763;
          lut[2978] <= 16'd15991;
          lut[2979] <= 16'd16211;
          lut[2980] <= 16'd16421;
          lut[2981] <= 16'd16624;
          lut[2982] <= 16'd16818;
          lut[2983] <= 16'd17006;
          lut[2984] <= 16'd17186;
          lut[2985] <= 16'd17360;
          lut[2986] <= 16'd17527;
          lut[2987] <= 16'd17689;
          lut[2988] <= 16'd17844;
          lut[2989] <= 16'd17995;
          lut[2990] <= 16'd18140;
          lut[2991] <= 16'd18280;
          lut[2992] <= 16'd18415;
          lut[2993] <= 16'd18546;
          lut[2994] <= 16'd18672;
          lut[2995] <= 16'd18795;
          lut[2996] <= 16'd18913;
          lut[2997] <= 16'd19028;
          lut[2998] <= 16'd19139;
          lut[2999] <= 16'd19247;
          lut[3000] <= 16'd19351;
          lut[3001] <= 16'd19452;
          lut[3002] <= 16'd19550;
          lut[3003] <= 16'd19646;
          lut[3004] <= 16'd19738;
          lut[3005] <= 16'd19828;
          lut[3006] <= 16'd19916;
          lut[3007] <= 16'd20001;
          lut[3008] <= 16'd20083;
          lut[3009] <= 16'd20164;
          lut[3010] <= 16'd20242;
          lut[3011] <= 16'd20318;
          lut[3012] <= 16'd20392;
          lut[3013] <= 16'd20464;
          lut[3014] <= 16'd20535;
          lut[3015] <= 16'd20603;
          lut[3016] <= 16'd20670;
          lut[3017] <= 16'd20735;
          lut[3018] <= 16'd20799;
          lut[3019] <= 16'd20861;
          lut[3020] <= 16'd20921;
          lut[3021] <= 16'd20980;
          lut[3022] <= 16'd21038;
          lut[3023] <= 16'd21094;
          lut[3024] <= 16'd21149;
          lut[3025] <= 16'd21203;
          lut[3026] <= 16'd21256;
          lut[3027] <= 16'd21307;
          lut[3028] <= 16'd21357;
          lut[3029] <= 16'd21406;
          lut[3030] <= 16'd21454;
          lut[3031] <= 16'd21501;
          lut[3032] <= 16'd21547;
          lut[3033] <= 16'd21593;
          lut[3034] <= 16'd21637;
          lut[3035] <= 16'd21680;
          lut[3036] <= 16'd21722;
          lut[3037] <= 16'd21764;
          lut[3038] <= 16'd21804;
          lut[3039] <= 16'd21844;
          lut[3040] <= 16'd21883;
          lut[3041] <= 16'd21922;
          lut[3042] <= 16'd21959;
          lut[3043] <= 16'd21996;
          lut[3044] <= 16'd22032;
          lut[3045] <= 16'd22067;
          lut[3046] <= 16'd22102;
          lut[3047] <= 16'd22136;
          lut[3048] <= 16'd22170;
          lut[3049] <= 16'd22203;
          lut[3050] <= 16'd22235;
          lut[3051] <= 16'd22267;
          lut[3052] <= 16'd22298;
          lut[3053] <= 16'd22329;
          lut[3054] <= 16'd22359;
          lut[3055] <= 16'd22388;
          lut[3056] <= 16'd22417;
          lut[3057] <= 16'd22446;
          lut[3058] <= 16'd22474;
          lut[3059] <= 16'd22502;
          lut[3060] <= 16'd22529;
          lut[3061] <= 16'd22556;
          lut[3062] <= 16'd22582;
          lut[3063] <= 16'd22608;
          lut[3064] <= 16'd22633;
          lut[3065] <= 16'd22658;
          lut[3066] <= 16'd22683;
          lut[3067] <= 16'd22707;
          lut[3068] <= 16'd22731;
          lut[3069] <= 16'd22755;
          lut[3070] <= 16'd22778;
          lut[3071] <= 16'd22801;
          lut[3072] <= 0;
          lut[3073] <= 16'd682;
          lut[3074] <= 16'd1362;
          lut[3075] <= 16'd2037;
          lut[3076] <= 16'd2706;
          lut[3077] <= 16'd3365;
          lut[3078] <= 16'd4014;
          lut[3079] <= 16'd4650;
          lut[3080] <= 16'd5272;
          lut[3081] <= 16'd5878;
          lut[3082] <= 16'd6468;
          lut[3083] <= 16'd7041;
          lut[3084] <= 16'd7596;
          lut[3085] <= 16'd8133;
          lut[3086] <= 16'd8652;
          lut[3087] <= 16'd9152;
          lut[3088] <= 16'd9634;
          lut[3089] <= 16'd10097;
          lut[3090] <= 16'd10543;
          lut[3091] <= 16'd10971;
          lut[3092] <= 16'd11383;
          lut[3093] <= 16'd11777;
          lut[3094] <= 16'd12156;
          lut[3095] <= 16'd12519;
          lut[3096] <= 16'd12868;
          lut[3097] <= 16'd13202;
          lut[3098] <= 16'd13523;
          lut[3099] <= 16'd13831;
          lut[3100] <= 16'd14126;
          lut[3101] <= 16'd14409;
          lut[3102] <= 16'd14681;
          lut[3103] <= 16'd14942;
          lut[3104] <= 16'd15193;
          lut[3105] <= 16'd15434;
          lut[3106] <= 16'd15665;
          lut[3107] <= 16'd15888;
          lut[3108] <= 16'd16102;
          lut[3109] <= 16'd16308;
          lut[3110] <= 16'd16507;
          lut[3111] <= 16'd16698;
          lut[3112] <= 16'd16882;
          lut[3113] <= 16'd17059;
          lut[3114] <= 16'd17230;
          lut[3115] <= 16'd17395;
          lut[3116] <= 16'd17555;
          lut[3117] <= 16'd17708;
          lut[3118] <= 16'd17857;
          lut[3119] <= 16'd18001;
          lut[3120] <= 16'd18140;
          lut[3121] <= 16'd18274;
          lut[3122] <= 16'd18404;
          lut[3123] <= 16'd18530;
          lut[3124] <= 16'd18651;
          lut[3125] <= 16'd18769;
          lut[3126] <= 16'd18884;
          lut[3127] <= 16'd18995;
          lut[3128] <= 16'd19102;
          lut[3129] <= 16'd19207;
          lut[3130] <= 16'd19308;
          lut[3131] <= 16'd19406;
          lut[3132] <= 16'd19502;
          lut[3133] <= 16'd19595;
          lut[3134] <= 16'd19685;
          lut[3135] <= 16'd19772;
          lut[3136] <= 16'd19858;
          lut[3137] <= 16'd19941;
          lut[3138] <= 16'd20022;
          lut[3139] <= 16'd20100;
          lut[3140] <= 16'd20177;
          lut[3141] <= 16'd20252;
          lut[3142] <= 16'd20324;
          lut[3143] <= 16'd20395;
          lut[3144] <= 16'd20464;
          lut[3145] <= 16'd20532;
          lut[3146] <= 16'd20598;
          lut[3147] <= 16'd20662;
          lut[3148] <= 16'd20724;
          lut[3149] <= 16'd20786;
          lut[3150] <= 16'd20845;
          lut[3151] <= 16'd20904;
          lut[3152] <= 16'd20961;
          lut[3153] <= 16'd21016;
          lut[3154] <= 16'd21071;
          lut[3155] <= 16'd21124;
          lut[3156] <= 16'd21176;
          lut[3157] <= 16'd21227;
          lut[3158] <= 16'd21277;
          lut[3159] <= 16'd21326;
          lut[3160] <= 16'd21374;
          lut[3161] <= 16'd21420;
          lut[3162] <= 16'd21466;
          lut[3163] <= 16'd21511;
          lut[3164] <= 16'd21555;
          lut[3165] <= 16'd21598;
          lut[3166] <= 16'd21640;
          lut[3167] <= 16'd21682;
          lut[3168] <= 16'd21722;
          lut[3169] <= 16'd21762;
          lut[3170] <= 16'd21801;
          lut[3171] <= 16'd21839;
          lut[3172] <= 16'd21877;
          lut[3173] <= 16'd21914;
          lut[3174] <= 16'd21950;
          lut[3175] <= 16'd21985;
          lut[3176] <= 16'd22020;
          lut[3177] <= 16'd22054;
          lut[3178] <= 16'd22088;
          lut[3179] <= 16'd22121;
          lut[3180] <= 16'd22153;
          lut[3181] <= 16'd22185;
          lut[3182] <= 16'd22216;
          lut[3183] <= 16'd22247;
          lut[3184] <= 16'd22277;
          lut[3185] <= 16'd22307;
          lut[3186] <= 16'd22336;
          lut[3187] <= 16'd22365;
          lut[3188] <= 16'd22393;
          lut[3189] <= 16'd22421;
          lut[3190] <= 16'd22448;
          lut[3191] <= 16'd22475;
          lut[3192] <= 16'd22502;
          lut[3193] <= 16'd22528;
          lut[3194] <= 16'd22553;
          lut[3195] <= 16'd22579;
          lut[3196] <= 16'd22604;
          lut[3197] <= 16'd22628;
          lut[3198] <= 16'd22652;
          lut[3199] <= 16'd22676;
          lut[3200] <= 0;
          lut[3201] <= 16'd655;
          lut[3202] <= 16'd1308;
          lut[3203] <= 16'd1957;
          lut[3204] <= 16'd2599;
          lut[3205] <= 16'd3234;
          lut[3206] <= 16'd3859;
          lut[3207] <= 16'd4473;
          lut[3208] <= 16'd5074;
          lut[3209] <= 16'd5662;
          lut[3210] <= 16'd6234;
          lut[3211] <= 16'd6791;
          lut[3212] <= 16'd7332;
          lut[3213] <= 16'd7856;
          lut[3214] <= 16'd8364;
          lut[3215] <= 16'd8854;
          lut[3216] <= 16'd9328;
          lut[3217] <= 16'd9784;
          lut[3218] <= 16'd10224;
          lut[3219] <= 16'd10647;
          lut[3220] <= 16'd11055;
          lut[3221] <= 16'd11447;
          lut[3222] <= 16'd11824;
          lut[3223] <= 16'd12186;
          lut[3224] <= 16'd12534;
          lut[3225] <= 16'd12868;
          lut[3226] <= 16'd13189;
          lut[3227] <= 16'd13498;
          lut[3228] <= 16'd13794;
          lut[3229] <= 16'd14079;
          lut[3230] <= 16'd14353;
          lut[3231] <= 16'd14617;
          lut[3232] <= 16'd14870;
          lut[3233] <= 16'd15114;
          lut[3234] <= 16'd15348;
          lut[3235] <= 16'd15574;
          lut[3236] <= 16'd15791;
          lut[3237] <= 16'd16000;
          lut[3238] <= 16'd16202;
          lut[3239] <= 16'd16396;
          lut[3240] <= 16'd16584;
          lut[3241] <= 16'd16765;
          lut[3242] <= 16'd16939;
          lut[3243] <= 16'd17108;
          lut[3244] <= 16'd17270;
          lut[3245] <= 16'd17428;
          lut[3246] <= 16'd17580;
          lut[3247] <= 16'd17727;
          lut[3248] <= 16'd17869;
          lut[3249] <= 16'd18006;
          lut[3250] <= 16'd18140;
          lut[3251] <= 16'd18269;
          lut[3252] <= 16'd18394;
          lut[3253] <= 16'd18515;
          lut[3254] <= 16'd18632;
          lut[3255] <= 16'd18746;
          lut[3256] <= 16'd18857;
          lut[3257] <= 16'd18964;
          lut[3258] <= 16'd19068;
          lut[3259] <= 16'd19169;
          lut[3260] <= 16'd19268;
          lut[3261] <= 16'd19363;
          lut[3262] <= 16'd19456;
          lut[3263] <= 16'd19547;
          lut[3264] <= 16'd19635;
          lut[3265] <= 16'd19720;
          lut[3266] <= 16'd19803;
          lut[3267] <= 16'd19885;
          lut[3268] <= 16'd19964;
          lut[3269] <= 16'd20041;
          lut[3270] <= 16'd20116;
          lut[3271] <= 16'd20189;
          lut[3272] <= 16'd20260;
          lut[3273] <= 16'd20330;
          lut[3274] <= 16'd20398;
          lut[3275] <= 16'd20464;
          lut[3276] <= 16'd20529;
          lut[3277] <= 16'd20592;
          lut[3278] <= 16'd20654;
          lut[3279] <= 16'd20714;
          lut[3280] <= 16'd20773;
          lut[3281] <= 16'd20831;
          lut[3282] <= 16'd20887;
          lut[3283] <= 16'd20943;
          lut[3284] <= 16'd20997;
          lut[3285] <= 16'd21049;
          lut[3286] <= 16'd21101;
          lut[3287] <= 16'd21151;
          lut[3288] <= 16'd21201;
          lut[3289] <= 16'd21249;
          lut[3290] <= 16'd21297;
          lut[3291] <= 16'd21343;
          lut[3292] <= 16'd21389;
          lut[3293] <= 16'd21433;
          lut[3294] <= 16'd21477;
          lut[3295] <= 16'd21520;
          lut[3296] <= 16'd21562;
          lut[3297] <= 16'd21603;
          lut[3298] <= 16'd21644;
          lut[3299] <= 16'd21683;
          lut[3300] <= 16'd21722;
          lut[3301] <= 16'd21760;
          lut[3302] <= 16'd21798;
          lut[3303] <= 16'd21835;
          lut[3304] <= 16'd21871;
          lut[3305] <= 16'd21906;
          lut[3306] <= 16'd21941;
          lut[3307] <= 16'd21975;
          lut[3308] <= 16'd22009;
          lut[3309] <= 16'd22042;
          lut[3310] <= 16'd22074;
          lut[3311] <= 16'd22106;
          lut[3312] <= 16'd22138;
          lut[3313] <= 16'd22169;
          lut[3314] <= 16'd22199;
          lut[3315] <= 16'd22229;
          lut[3316] <= 16'd22258;
          lut[3317] <= 16'd22287;
          lut[3318] <= 16'd22315;
          lut[3319] <= 16'd22343;
          lut[3320] <= 16'd22371;
          lut[3321] <= 16'd22398;
          lut[3322] <= 16'd22424;
          lut[3323] <= 16'd22451;
          lut[3324] <= 16'd22476;
          lut[3325] <= 16'd22502;
          lut[3326] <= 16'd22527;
          lut[3327] <= 16'd22551;
          lut[3328] <= 0;
          lut[3329] <= 16'd630;
          lut[3330] <= 16'd1258;
          lut[3331] <= 16'd1882;
          lut[3332] <= 16'd2501;
          lut[3333] <= 16'd3113;
          lut[3334] <= 16'd3716;
          lut[3335] <= 16'd4309;
          lut[3336] <= 16'd4891;
          lut[3337] <= 16'd5460;
          lut[3338] <= 16'd6016;
          lut[3339] <= 16'd6558;
          lut[3340] <= 16'd7085;
          lut[3341] <= 16'd7596;
          lut[3342] <= 16'd8093;
          lut[3343] <= 16'd8573;
          lut[3344] <= 16'd9038;
          lut[3345] <= 16'd9488;
          lut[3346] <= 16'd9921;
          lut[3347] <= 16'd10340;
          lut[3348] <= 16'd10743;
          lut[3349] <= 16'd11132;
          lut[3350] <= 16'd11506;
          lut[3351] <= 16'd11866;
          lut[3352] <= 16'd12213;
          lut[3353] <= 16'd12547;
          lut[3354] <= 16'd12868;
          lut[3355] <= 16'd13177;
          lut[3356] <= 16'd13475;
          lut[3357] <= 16'd13761;
          lut[3358] <= 16'd14036;
          lut[3359] <= 16'd14301;
          lut[3360] <= 16'd14557;
          lut[3361] <= 16'd14803;
          lut[3362] <= 16'd15040;
          lut[3363] <= 16'd15268;
          lut[3364] <= 16'd15488;
          lut[3365] <= 16'd15700;
          lut[3366] <= 16'd15905;
          lut[3367] <= 16'd16102;
          lut[3368] <= 16'd16293;
          lut[3369] <= 16'd16477;
          lut[3370] <= 16'd16654;
          lut[3371] <= 16'd16826;
          lut[3372] <= 16'd16992;
          lut[3373] <= 16'd17152;
          lut[3374] <= 16'd17307;
          lut[3375] <= 16'd17457;
          lut[3376] <= 16'd17603;
          lut[3377] <= 16'd17743;
          lut[3378] <= 16'd17879;
          lut[3379] <= 16'd18012;
          lut[3380] <= 16'd18140;
          lut[3381] <= 16'd18264;
          lut[3382] <= 16'd18384;
          lut[3383] <= 16'd18501;
          lut[3384] <= 16'd18614;
          lut[3385] <= 16'd18724;
          lut[3386] <= 16'd18831;
          lut[3387] <= 16'd18935;
          lut[3388] <= 16'd19036;
          lut[3389] <= 16'd19135;
          lut[3390] <= 16'd19230;
          lut[3391] <= 16'd19323;
          lut[3392] <= 16'd19414;
          lut[3393] <= 16'd19502;
          lut[3394] <= 16'd19587;
          lut[3395] <= 16'd19671;
          lut[3396] <= 16'd19752;
          lut[3397] <= 16'd19832;
          lut[3398] <= 16'd19909;
          lut[3399] <= 16'd19985;
          lut[3400] <= 16'd20058;
          lut[3401] <= 16'd20130;
          lut[3402] <= 16'd20200;
          lut[3403] <= 16'd20269;
          lut[3404] <= 16'd20335;
          lut[3405] <= 16'd20401;
          lut[3406] <= 16'd20464;
          lut[3407] <= 16'd20527;
          lut[3408] <= 16'd20588;
          lut[3409] <= 16'd20647;
          lut[3410] <= 16'd20705;
          lut[3411] <= 16'd20762;
          lut[3412] <= 16'd20818;
          lut[3413] <= 16'd20872;
          lut[3414] <= 16'd20926;
          lut[3415] <= 16'd20978;
          lut[3416] <= 16'd21029;
          lut[3417] <= 16'd21079;
          lut[3418] <= 16'd21128;
          lut[3419] <= 16'd21176;
          lut[3420] <= 16'd21223;
          lut[3421] <= 16'd21269;
          lut[3422] <= 16'd21315;
          lut[3423] <= 16'd21359;
          lut[3424] <= 16'd21403;
          lut[3425] <= 16'd21445;
          lut[3426] <= 16'd21487;
          lut[3427] <= 16'd21528;
          lut[3428] <= 16'd21568;
          lut[3429] <= 16'd21608;
          lut[3430] <= 16'd21647;
          lut[3431] <= 16'd21685;
          lut[3432] <= 16'd21722;
          lut[3433] <= 16'd21759;
          lut[3434] <= 16'd21795;
          lut[3435] <= 16'd21830;
          lut[3436] <= 16'd21865;
          lut[3437] <= 16'd21900;
          lut[3438] <= 16'd21933;
          lut[3439] <= 16'd21966;
          lut[3440] <= 16'd21999;
          lut[3441] <= 16'd22031;
          lut[3442] <= 16'd22062;
          lut[3443] <= 16'd22093;
          lut[3444] <= 16'd22123;
          lut[3445] <= 16'd22153;
          lut[3446] <= 16'd22183;
          lut[3447] <= 16'd22212;
          lut[3448] <= 16'd22240;
          lut[3449] <= 16'd22268;
          lut[3450] <= 16'd22296;
          lut[3451] <= 16'd22323;
          lut[3452] <= 16'd22350;
          lut[3453] <= 16'd22376;
          lut[3454] <= 16'd22402;
          lut[3455] <= 16'd22427;
          lut[3456] <= 0;
          lut[3457] <= 16'd607;
          lut[3458] <= 16'd1211;
          lut[3459] <= 16'd1813;
          lut[3460] <= 16'd2410;
          lut[3461] <= 16'd3000;
          lut[3462] <= 16'd3583;
          lut[3463] <= 16'd4156;
          lut[3464] <= 16'd4720;
          lut[3465] <= 16'd5272;
          lut[3466] <= 16'd5811;
          lut[3467] <= 16'd6339;
          lut[3468] <= 16'd6852;
          lut[3469] <= 16'd7352;
          lut[3470] <= 16'd7837;
          lut[3471] <= 16'd8308;
          lut[3472] <= 16'd8765;
          lut[3473] <= 16'd9207;
          lut[3474] <= 16'd9634;
          lut[3475] <= 16'd10047;
          lut[3476] <= 16'd10446;
          lut[3477] <= 16'd10831;
          lut[3478] <= 16'd11202;
          lut[3479] <= 16'd11560;
          lut[3480] <= 16'd11905;
          lut[3481] <= 16'd12238;
          lut[3482] <= 16'd12559;
          lut[3483] <= 16'd12868;
          lut[3484] <= 16'd13166;
          lut[3485] <= 16'd13453;
          lut[3486] <= 16'd13729;
          lut[3487] <= 16'd13996;
          lut[3488] <= 16'd14253;
          lut[3489] <= 16'd14501;
          lut[3490] <= 16'd14740;
          lut[3491] <= 16'd14970;
          lut[3492] <= 16'd15193;
          lut[3493] <= 16'd15407;
          lut[3494] <= 16'd15615;
          lut[3495] <= 16'd15815;
          lut[3496] <= 16'd16008;
          lut[3497] <= 16'd16195;
          lut[3498] <= 16'd16375;
          lut[3499] <= 16'd16550;
          lut[3500] <= 16'd16718;
          lut[3501] <= 16'd16882;
          lut[3502] <= 16'd17040;
          lut[3503] <= 16'd17193;
          lut[3504] <= 16'd17341;
          lut[3505] <= 16'd17485;
          lut[3506] <= 16'd17624;
          lut[3507] <= 16'd17759;
          lut[3508] <= 16'd17889;
          lut[3509] <= 16'd18016;
          lut[3510] <= 16'd18140;
          lut[3511] <= 16'd18259;
          lut[3512] <= 16'd18375;
          lut[3513] <= 16'd18488;
          lut[3514] <= 16'd18598;
          lut[3515] <= 16'd18704;
          lut[3516] <= 16'd18808;
          lut[3517] <= 16'd18909;
          lut[3518] <= 16'd19007;
          lut[3519] <= 16'd19102;
          lut[3520] <= 16'd19195;
          lut[3521] <= 16'd19286;
          lut[3522] <= 16'd19374;
          lut[3523] <= 16'd19460;
          lut[3524] <= 16'd19543;
          lut[3525] <= 16'd19625;
          lut[3526] <= 16'd19704;
          lut[3527] <= 16'd19782;
          lut[3528] <= 16'd19858;
          lut[3529] <= 16'd19932;
          lut[3530] <= 16'd20004;
          lut[3531] <= 16'd20074;
          lut[3532] <= 16'd20143;
          lut[3533] <= 16'd20210;
          lut[3534] <= 16'd20276;
          lut[3535] <= 16'd20340;
          lut[3536] <= 16'd20403;
          lut[3537] <= 16'd20464;
          lut[3538] <= 16'd20524;
          lut[3539] <= 16'd20583;
          lut[3540] <= 16'd20641;
          lut[3541] <= 16'd20697;
          lut[3542] <= 16'd20752;
          lut[3543] <= 16'd20806;
          lut[3544] <= 16'd20858;
          lut[3545] <= 16'd20910;
          lut[3546] <= 16'd20961;
          lut[3547] <= 16'd21010;
          lut[3548] <= 16'd21059;
          lut[3549] <= 16'd21107;
          lut[3550] <= 16'd21153;
          lut[3551] <= 16'd21199;
          lut[3552] <= 16'd21244;
          lut[3553] <= 16'd21288;
          lut[3554] <= 16'd21331;
          lut[3555] <= 16'd21374;
          lut[3556] <= 16'd21415;
          lut[3557] <= 16'd21456;
          lut[3558] <= 16'd21496;
          lut[3559] <= 16'd21536;
          lut[3560] <= 16'd21574;
          lut[3561] <= 16'd21612;
          lut[3562] <= 16'd21650;
          lut[3563] <= 16'd21686;
          lut[3564] <= 16'd21722;
          lut[3565] <= 16'd21758;
          lut[3566] <= 16'd21792;
          lut[3567] <= 16'd21827;
          lut[3568] <= 16'd21860;
          lut[3569] <= 16'd21893;
          lut[3570] <= 16'd21926;
          lut[3571] <= 16'd21958;
          lut[3572] <= 16'd21989;
          lut[3573] <= 16'd22020;
          lut[3574] <= 16'd22050;
          lut[3575] <= 16'd22080;
          lut[3576] <= 16'd22110;
          lut[3577] <= 16'd22139;
          lut[3578] <= 16'd22167;
          lut[3579] <= 16'd22196;
          lut[3580] <= 16'd22223;
          lut[3581] <= 16'd22251;
          lut[3582] <= 16'd22277;
          lut[3583] <= 16'd22304;
          lut[3584] <= 0;
          lut[3585] <= 16'd585;
          lut[3586] <= 16'd1168;
          lut[3587] <= 16'd1749;
          lut[3588] <= 16'd2325;
          lut[3589] <= 16'd2895;
          lut[3590] <= 16'd3459;
          lut[3591] <= 16'd4014;
          lut[3592] <= 16'd4560;
          lut[3593] <= 16'd5095;
          lut[3594] <= 16'd5620;
          lut[3595] <= 16'd6133;
          lut[3596] <= 16'd6634;
          lut[3597] <= 16'd7122;
          lut[3598] <= 16'd7596;
          lut[3599] <= 16'd8058;
          lut[3600] <= 16'd8506;
          lut[3601] <= 16'd8940;
          lut[3602] <= 16'd9361;
          lut[3603] <= 16'd9768;
          lut[3604] <= 16'd10162;
          lut[3605] <= 16'd10543;
          lut[3606] <= 16'd10911;
          lut[3607] <= 16'd11267;
          lut[3608] <= 16'd11610;
          lut[3609] <= 16'd11942;
          lut[3610] <= 16'd12261;
          lut[3611] <= 16'd12570;
          lut[3612] <= 16'd12868;
          lut[3613] <= 16'd13155;
          lut[3614] <= 16'd13433;
          lut[3615] <= 16'd13700;
          lut[3616] <= 16'd13959;
          lut[3617] <= 16'd14208;
          lut[3618] <= 16'd14449;
          lut[3619] <= 16'd14681;
          lut[3620] <= 16'd14905;
          lut[3621] <= 16'd15122;
          lut[3622] <= 16'd15332;
          lut[3623] <= 16'd15534;
          lut[3624] <= 16'd15730;
          lut[3625] <= 16'd15919;
          lut[3626] <= 16'd16102;
          lut[3627] <= 16'd16279;
          lut[3628] <= 16'd16451;
          lut[3629] <= 16'd16617;
          lut[3630] <= 16'd16777;
          lut[3631] <= 16'd16933;
          lut[3632] <= 16'd17084;
          lut[3633] <= 16'd17230;
          lut[3634] <= 16'd17372;
          lut[3635] <= 16'd17510;
          lut[3636] <= 16'd17643;
          lut[3637] <= 16'd17773;
          lut[3638] <= 16'd17899;
          lut[3639] <= 16'd18021;
          lut[3640] <= 16'd18140;
          lut[3641] <= 16'd18255;
          lut[3642] <= 16'd18367;
          lut[3643] <= 16'd18476;
          lut[3644] <= 16'd18582;
          lut[3645] <= 16'd18685;
          lut[3646] <= 16'd18786;
          lut[3647] <= 16'd18884;
          lut[3648] <= 16'd18979;
          lut[3649] <= 16'd19072;
          lut[3650] <= 16'd19162;
          lut[3651] <= 16'd19250;
          lut[3652] <= 16'd19336;
          lut[3653] <= 16'd19420;
          lut[3654] <= 16'd19502;
          lut[3655] <= 16'd19581;
          lut[3656] <= 16'd19659;
          lut[3657] <= 16'd19735;
          lut[3658] <= 16'd19809;
          lut[3659] <= 16'd19882;
          lut[3660] <= 16'd19953;
          lut[3661] <= 16'd20022;
          lut[3662] <= 16'd20089;
          lut[3663] <= 16'd20155;
          lut[3664] <= 16'd20220;
          lut[3665] <= 16'd20283;
          lut[3666] <= 16'd20345;
          lut[3667] <= 16'd20405;
          lut[3668] <= 16'd20464;
          lut[3669] <= 16'd20522;
          lut[3670] <= 16'd20579;
          lut[3671] <= 16'd20634;
          lut[3672] <= 16'd20689;
          lut[3673] <= 16'd20742;
          lut[3674] <= 16'd20794;
          lut[3675] <= 16'd20845;
          lut[3676] <= 16'd20895;
          lut[3677] <= 16'd20945;
          lut[3678] <= 16'd20993;
          lut[3679] <= 16'd21040;
          lut[3680] <= 16'd21086;
          lut[3681] <= 16'd21132;
          lut[3682] <= 16'd21176;
          lut[3683] <= 16'd21220;
          lut[3684] <= 16'd21263;
          lut[3685] <= 16'd21305;
          lut[3686] <= 16'd21346;
          lut[3687] <= 16'd21387;
          lut[3688] <= 16'd21427;
          lut[3689] <= 16'd21466;
          lut[3690] <= 16'd21505;
          lut[3691] <= 16'd21543;
          lut[3692] <= 16'd21580;
          lut[3693] <= 16'd21616;
          lut[3694] <= 16'd21652;
          lut[3695] <= 16'd21687;
          lut[3696] <= 16'd21722;
          lut[3697] <= 16'd21756;
          lut[3698] <= 16'd21790;
          lut[3699] <= 16'd21823;
          lut[3700] <= 16'd21855;
          lut[3701] <= 16'd21887;
          lut[3702] <= 16'd21919;
          lut[3703] <= 16'd21950;
          lut[3704] <= 16'd21980;
          lut[3705] <= 16'd22010;
          lut[3706] <= 16'd22040;
          lut[3707] <= 16'd22069;
          lut[3708] <= 16'd22097;
          lut[3709] <= 16'd22126;
          lut[3710] <= 16'd22153;
          lut[3711] <= 16'd22181;
          lut[3712] <= 0;
          lut[3713] <= 16'd565;
          lut[3714] <= 16'd1128;
          lut[3715] <= 16'd1689;
          lut[3716] <= 16'd2246;
          lut[3717] <= 16'd2797;
          lut[3718] <= 16'd3343;
          lut[3719] <= 16'd3881;
          lut[3720] <= 16'd4410;
          lut[3721] <= 16'd4930;
          lut[3722] <= 16'd5440;
          lut[3723] <= 16'd5940;
          lut[3724] <= 16'd6428;
          lut[3725] <= 16'd6905;
          lut[3726] <= 16'd7369;
          lut[3727] <= 16'd7821;
          lut[3728] <= 16'd8260;
          lut[3729] <= 16'd8687;
          lut[3730] <= 16'd9101;
          lut[3731] <= 16'd9503;
          lut[3732] <= 16'd9892;
          lut[3733] <= 16'd10269;
          lut[3734] <= 16'd10633;
          lut[3735] <= 16'd10986;
          lut[3736] <= 16'd11327;
          lut[3737] <= 16'd11657;
          lut[3738] <= 16'd11975;
          lut[3739] <= 16'd12283;
          lut[3740] <= 16'd12581;
          lut[3741] <= 16'd12868;
          lut[3742] <= 16'd13146;
          lut[3743] <= 16'd13414;
          lut[3744] <= 16'd13673;
          lut[3745] <= 16'd13924;
          lut[3746] <= 16'd14166;
          lut[3747] <= 16'd14399;
          lut[3748] <= 16'd14626;
          lut[3749] <= 16'd14844;
          lut[3750] <= 16'd15056;
          lut[3751] <= 16'd15260;
          lut[3752] <= 16'd15458;
          lut[3753] <= 16'd15650;
          lut[3754] <= 16'd15835;
          lut[3755] <= 16'd16014;
          lut[3756] <= 16'd16188;
          lut[3757] <= 16'd16357;
          lut[3758] <= 16'd16520;
          lut[3759] <= 16'd16678;
          lut[3760] <= 16'd16832;
          lut[3761] <= 16'd16980;
          lut[3762] <= 16'd17125;
          lut[3763] <= 16'd17265;
          lut[3764] <= 16'd17401;
          lut[3765] <= 16'd17533;
          lut[3766] <= 16'd17661;
          lut[3767] <= 16'd17786;
          lut[3768] <= 16'd17907;
          lut[3769] <= 16'd18025;
          lut[3770] <= 16'd18140;
          lut[3771] <= 16'd18251;
          lut[3772] <= 16'd18359;
          lut[3773] <= 16'd18465;
          lut[3774] <= 16'd18568;
          lut[3775] <= 16'd18668;
          lut[3776] <= 16'd18765;
          lut[3777] <= 16'd18860;
          lut[3778] <= 16'd18953;
          lut[3779] <= 16'd19043;
          lut[3780] <= 16'd19131;
          lut[3781] <= 16'd19217;
          lut[3782] <= 16'd19301;
          lut[3783] <= 16'd19383;
          lut[3784] <= 16'd19463;
          lut[3785] <= 16'd19540;
          lut[3786] <= 16'd19617;
          lut[3787] <= 16'd19691;
          lut[3788] <= 16'd19764;
          lut[3789] <= 16'd19835;
          lut[3790] <= 16'd19904;
          lut[3791] <= 16'd19972;
          lut[3792] <= 16'd20038;
          lut[3793] <= 16'd20103;
          lut[3794] <= 16'd20167;
          lut[3795] <= 16'd20229;
          lut[3796] <= 16'd20289;
          lut[3797] <= 16'd20349;
          lut[3798] <= 16'd20407;
          lut[3799] <= 16'd20464;
          lut[3800] <= 16'd20520;
          lut[3801] <= 16'd20575;
          lut[3802] <= 16'd20629;
          lut[3803] <= 16'd20681;
          lut[3804] <= 16'd20733;
          lut[3805] <= 16'd20783;
          lut[3806] <= 16'd20833;
          lut[3807] <= 16'd20882;
          lut[3808] <= 16'd20929;
          lut[3809] <= 16'd20976;
          lut[3810] <= 16'd21022;
          lut[3811] <= 16'd21067;
          lut[3812] <= 16'd21111;
          lut[3813] <= 16'd21155;
          lut[3814] <= 16'd21197;
          lut[3815] <= 16'd21239;
          lut[3816] <= 16'd21280;
          lut[3817] <= 16'd21321;
          lut[3818] <= 16'd21361;
          lut[3819] <= 16'd21400;
          lut[3820] <= 16'd21438;
          lut[3821] <= 16'd21476;
          lut[3822] <= 16'd21513;
          lut[3823] <= 16'd21549;
          lut[3824] <= 16'd21585;
          lut[3825] <= 16'd21620;
          lut[3826] <= 16'd21655;
          lut[3827] <= 16'd21689;
          lut[3828] <= 16'd21722;
          lut[3829] <= 16'd21755;
          lut[3830] <= 16'd21788;
          lut[3831] <= 16'd21820;
          lut[3832] <= 16'd21851;
          lut[3833] <= 16'd21882;
          lut[3834] <= 16'd21912;
          lut[3835] <= 16'd21942;
          lut[3836] <= 16'd21972;
          lut[3837] <= 16'd22001;
          lut[3838] <= 16'd22030;
          lut[3839] <= 16'd22058;
          lut[3840] <= 0;
          lut[3841] <= 16'd546;
          lut[3842] <= 16'd1091;
          lut[3843] <= 16'd1633;
          lut[3844] <= 16'd2172;
          lut[3845] <= 16'd2706;
          lut[3846] <= 16'd3234;
          lut[3847] <= 16'd3756;
          lut[3848] <= 16'd4270;
          lut[3849] <= 16'd4775;
          lut[3850] <= 16'd5272;
          lut[3851] <= 16'd5758;
          lut[3852] <= 16'd6234;
          lut[3853] <= 16'd6700;
          lut[3854] <= 16'd7154;
          lut[3855] <= 16'd7596;
          lut[3856] <= 16'd8027;
          lut[3857] <= 16'd8447;
          lut[3858] <= 16'd8854;
          lut[3859] <= 16'd9250;
          lut[3860] <= 16'd9634;
          lut[3861] <= 16'd10006;
          lut[3862] <= 16'd10367;
          lut[3863] <= 16'd10716;
          lut[3864] <= 16'd11055;
          lut[3865] <= 16'd11383;
          lut[3866] <= 16'd11700;
          lut[3867] <= 16'd12006;
          lut[3868] <= 16'd12303;
          lut[3869] <= 16'd12590;
          lut[3870] <= 16'd12868;
          lut[3871] <= 16'd13137;
          lut[3872] <= 16'd13396;
          lut[3873] <= 16'd13648;
          lut[3874] <= 16'd13891;
          lut[3875] <= 16'd14126;
          lut[3876] <= 16'd14353;
          lut[3877] <= 16'd14574;
          lut[3878] <= 16'd14787;
          lut[3879] <= 16'd14993;
          lut[3880] <= 16'd15193;
          lut[3881] <= 16'd15386;
          lut[3882] <= 16'd15574;
          lut[3883] <= 16'd15755;
          lut[3884] <= 16'd15931;
          lut[3885] <= 16'd16102;
          lut[3886] <= 16'd16268;
          lut[3887] <= 16'd16428;
          lut[3888] <= 16'd16584;
          lut[3889] <= 16'd16735;
          lut[3890] <= 16'd16882;
          lut[3891] <= 16'd17024;
          lut[3892] <= 16'd17163;
          lut[3893] <= 16'd17297;
          lut[3894] <= 16'd17428;
          lut[3895] <= 16'd17555;
          lut[3896] <= 16'd17678;
          lut[3897] <= 16'd17798;
          lut[3898] <= 16'd17915;
          lut[3899] <= 16'd18029;
          lut[3900] <= 16'd18140;
          lut[3901] <= 16'd18247;
          lut[3902] <= 16'd18352;
          lut[3903] <= 16'd18455;
          lut[3904] <= 16'd18554;
          lut[3905] <= 16'd18651;
          lut[3906] <= 16'd18746;
          lut[3907] <= 16'd18838;
          lut[3908] <= 16'd18929;
          lut[3909] <= 16'd19016;
          lut[3910] <= 16'd19102;
          lut[3911] <= 16'd19186;
          lut[3912] <= 16'd19268;
          lut[3913] <= 16'd19348;
          lut[3914] <= 16'd19426;
          lut[3915] <= 16'd19502;
          lut[3916] <= 16'd19576;
          lut[3917] <= 16'd19649;
          lut[3918] <= 16'd19720;
          lut[3919] <= 16'd19790;
          lut[3920] <= 16'd19858;
          lut[3921] <= 16'd19924;
          lut[3922] <= 16'd19990;
          lut[3923] <= 16'd20053;
          lut[3924] <= 16'd20116;
          lut[3925] <= 16'd20177;
          lut[3926] <= 16'd20237;
          lut[3927] <= 16'd20295;
          lut[3928] <= 16'd20353;
          lut[3929] <= 16'd20409;
          lut[3930] <= 16'd20464;
          lut[3931] <= 16'd20518;
          lut[3932] <= 16'd20571;
          lut[3933] <= 16'd20623;
          lut[3934] <= 16'd20674;
          lut[3935] <= 16'd20724;
          lut[3936] <= 16'd20773;
          lut[3937] <= 16'd20822;
          lut[3938] <= 16'd20869;
          lut[3939] <= 16'd20915;
          lut[3940] <= 16'd20961;
          lut[3941] <= 16'd21005;
          lut[3942] <= 16'd21049;
          lut[3943] <= 16'd21092;
          lut[3944] <= 16'd21135;
          lut[3945] <= 16'd21176;
          lut[3946] <= 16'd21217;
          lut[3947] <= 16'd21257;
          lut[3948] <= 16'd21297;
          lut[3949] <= 16'd21336;
          lut[3950] <= 16'd21374;
          lut[3951] <= 16'd21411;
          lut[3952] <= 16'd21448;
          lut[3953] <= 16'd21484;
          lut[3954] <= 16'd21520;
          lut[3955] <= 16'd21555;
          lut[3956] <= 16'd21590;
          lut[3957] <= 16'd21623;
          lut[3958] <= 16'd21657;
          lut[3959] <= 16'd21690;
          lut[3960] <= 16'd21722;
          lut[3961] <= 16'd21754;
          lut[3962] <= 16'd21785;
          lut[3963] <= 16'd21816;
          lut[3964] <= 16'd21847;
          lut[3965] <= 16'd21877;
          lut[3966] <= 16'd21906;
          lut[3967] <= 16'd21935;
          lut[3968] <= 0;
          lut[3969] <= 16'd528;
          lut[3970] <= 16'd1056;
          lut[3971] <= 16'd1581;
          lut[3972] <= 16'd2102;
          lut[3973] <= 16'd2620;
          lut[3974] <= 16'd3132;
          lut[3975] <= 16'd3639;
          lut[3976] <= 16'd4138;
          lut[3977] <= 16'd4629;
          lut[3978] <= 16'd5112;
          lut[3979] <= 16'd5587;
          lut[3980] <= 16'd6051;
          lut[3981] <= 16'd6506;
          lut[3982] <= 16'd6950;
          lut[3983] <= 16'd7384;
          lut[3984] <= 16'd7806;
          lut[3985] <= 16'd8218;
          lut[3986] <= 16'd8619;
          lut[3987] <= 16'd9009;
          lut[3988] <= 16'd9387;
          lut[3989] <= 16'd9755;
          lut[3990] <= 16'd10112;
          lut[3991] <= 16'd10458;
          lut[3992] <= 16'd10794;
          lut[3993] <= 16'd11119;
          lut[3994] <= 16'd11434;
          lut[3995] <= 16'd11740;
          lut[3996] <= 16'd12036;
          lut[3997] <= 16'd12322;
          lut[3998] <= 16'd12599;
          lut[3999] <= 16'd12868;
          lut[4000] <= 16'd13128;
          lut[4001] <= 16'd13380;
          lut[4002] <= 16'd13624;
          lut[4003] <= 16'd13860;
          lut[4004] <= 16'd14088;
          lut[4005] <= 16'd14310;
          lut[4006] <= 16'd14524;
          lut[4007] <= 16'd14732;
          lut[4008] <= 16'd14934;
          lut[4009] <= 16'd15129;
          lut[4010] <= 16'd15318;
          lut[4011] <= 16'd15502;
          lut[4012] <= 16'd15680;
          lut[4013] <= 16'd15853;
          lut[4014] <= 16'd16020;
          lut[4015] <= 16'd16183;
          lut[4016] <= 16'd16341;
          lut[4017] <= 16'd16494;
          lut[4018] <= 16'd16643;
          lut[4019] <= 16'd16788;
          lut[4020] <= 16'd16928;
          lut[4021] <= 16'd17065;
          lut[4022] <= 16'd17198;
          lut[4023] <= 16'd17327;
          lut[4024] <= 16'd17452;
          lut[4025] <= 16'd17575;
          lut[4026] <= 16'd17694;
          lut[4027] <= 16'd17810;
          lut[4028] <= 16'd17923;
          lut[4029] <= 16'd18032;
          lut[4030] <= 16'd18140;
          lut[4031] <= 16'd18244;
          lut[4032] <= 16'd18346;
          lut[4033] <= 16'd18445;
          lut[4034] <= 16'd18542;
          lut[4035] <= 16'd18636;
          lut[4036] <= 16'd18728;
          lut[4037] <= 16'd18818;
          lut[4038] <= 16'd18905;
          lut[4039] <= 16'd18991;
          lut[4040] <= 16'd19075;
          lut[4041] <= 16'd19156;
          lut[4042] <= 16'd19236;
          lut[4043] <= 16'd19314;
          lut[4044] <= 16'd19391;
          lut[4045] <= 16'd19465;
          lut[4046] <= 16'd19538;
          lut[4047] <= 16'd19609;
          lut[4048] <= 16'd19679;
          lut[4049] <= 16'd19747;
          lut[4050] <= 16'd19814;
          lut[4051] <= 16'd19879;
          lut[4052] <= 16'd19943;
          lut[4053] <= 16'd20006;
          lut[4054] <= 16'd20068;
          lut[4055] <= 16'd20128;
          lut[4056] <= 16'd20187;
          lut[4057] <= 16'd20244;
          lut[4058] <= 16'd20301;
          lut[4059] <= 16'd20357;
          lut[4060] <= 16'd20411;
          lut[4061] <= 16'd20464;
          lut[4062] <= 16'd20517;
          lut[4063] <= 16'd20568;
          lut[4064] <= 16'd20618;
          lut[4065] <= 16'd20668;
          lut[4066] <= 16'd20716;
          lut[4067] <= 16'd20764;
          lut[4068] <= 16'd20811;
          lut[4069] <= 16'd20857;
          lut[4070] <= 16'd20902;
          lut[4071] <= 16'd20946;
          lut[4072] <= 16'd20990;
          lut[4073] <= 16'd21032;
          lut[4074] <= 16'd21074;
          lut[4075] <= 16'd21116;
          lut[4076] <= 16'd21156;
          lut[4077] <= 16'd21196;
          lut[4078] <= 16'd21235;
          lut[4079] <= 16'd21274;
          lut[4080] <= 16'd21312;
          lut[4081] <= 16'd21349;
          lut[4082] <= 16'd21386;
          lut[4083] <= 16'd21422;
          lut[4084] <= 16'd21457;
          lut[4085] <= 16'd21492;
          lut[4086] <= 16'd21527;
          lut[4087] <= 16'd21561;
          lut[4088] <= 16'd21594;
          lut[4089] <= 16'd21627;
          lut[4090] <= 16'd21659;
          lut[4091] <= 16'd21691;
          lut[4092] <= 16'd21722;
          lut[4093] <= 16'd21753;
          lut[4094] <= 16'd21783;
          lut[4095] <= 16'd21813;
          lut[4096] <= 0;
          lut[4097] <= 16'd512;
          lut[4098] <= 16'd1023;
          lut[4099] <= 16'd1532;
          lut[4100] <= 16'd2037;
          lut[4101] <= 16'd2539;
          lut[4102] <= 16'd3037;
          lut[4103] <= 16'd3528;
          lut[4104] <= 16'd4014;
          lut[4105] <= 16'd4492;
          lut[4106] <= 16'd4962;
          lut[4107] <= 16'd5425;
          lut[4108] <= 16'd5878;
          lut[4109] <= 16'd6322;
          lut[4110] <= 16'd6757;
          lut[4111] <= 16'd7182;
          lut[4112] <= 16'd7596;
          lut[4113] <= 16'd8001;
          lut[4114] <= 16'd8395;
          lut[4115] <= 16'd8779;
          lut[4116] <= 16'd9152;
          lut[4117] <= 16'd9515;
          lut[4118] <= 16'd9868;
          lut[4119] <= 16'd10210;
          lut[4120] <= 16'd10543;
          lut[4121] <= 16'd10866;
          lut[4122] <= 16'd11179;
          lut[4123] <= 16'd11483;
          lut[4124] <= 16'd11777;
          lut[4125] <= 16'd12063;
          lut[4126] <= 16'd12340;
          lut[4127] <= 16'd12608;
          lut[4128] <= 16'd12868;
          lut[4129] <= 16'd13120;
          lut[4130] <= 16'd13364;
          lut[4131] <= 16'd13601;
          lut[4132] <= 16'd13831;
          lut[4133] <= 16'd14053;
          lut[4134] <= 16'd14269;
          lut[4135] <= 16'd14478;
          lut[4136] <= 16'd14681;
          lut[4137] <= 16'd14878;
          lut[4138] <= 16'd15069;
          lut[4139] <= 16'd15254;
          lut[4140] <= 16'd15434;
          lut[4141] <= 16'd15608;
          lut[4142] <= 16'd15778;
          lut[4143] <= 16'd15942;
          lut[4144] <= 16'd16102;
          lut[4145] <= 16'd16257;
          lut[4146] <= 16'd16408;
          lut[4147] <= 16'd16555;
          lut[4148] <= 16'd16698;
          lut[4149] <= 16'd16836;
          lut[4150] <= 16'd16971;
          lut[4151] <= 16'd17102;
          lut[4152] <= 16'd17230;
          lut[4153] <= 16'd17355;
          lut[4154] <= 16'd17476;
          lut[4155] <= 16'd17594;
          lut[4156] <= 16'd17708;
          lut[4157] <= 16'd17820;
          lut[4158] <= 16'd17929;
          lut[4159] <= 16'd18036;
          lut[4160] <= 16'd18140;
          lut[4161] <= 16'd18241;
          lut[4162] <= 16'd18339;
          lut[4163] <= 16'd18436;
          lut[4164] <= 16'd18530;
          lut[4165] <= 16'd18621;
          lut[4166] <= 16'd18711;
          lut[4167] <= 16'd18798;
          lut[4168] <= 16'd18884;
          lut[4169] <= 16'd18967;
          lut[4170] <= 16'd19049;
          lut[4171] <= 16'd19129;
          lut[4172] <= 16'd19207;
          lut[4173] <= 16'd19283;
          lut[4174] <= 16'd19357;
          lut[4175] <= 16'd19430;
          lut[4176] <= 16'd19502;
          lut[4177] <= 16'd19572;
          lut[4178] <= 16'd19640;
          lut[4179] <= 16'd19707;
          lut[4180] <= 16'd19772;
          lut[4181] <= 16'd19837;
          lut[4182] <= 16'd19900;
          lut[4183] <= 16'd19961;
          lut[4184] <= 16'd20022;
          lut[4185] <= 16'd20081;
          lut[4186] <= 16'd20139;
          lut[4187] <= 16'd20196;
          lut[4188] <= 16'd20252;
          lut[4189] <= 16'd20306;
          lut[4190] <= 16'd20360;
          lut[4191] <= 16'd20413;
          lut[4192] <= 16'd20464;
          lut[4193] <= 16'd20515;
          lut[4194] <= 16'd20565;
          lut[4195] <= 16'd20614;
          lut[4196] <= 16'd20662;
          lut[4197] <= 16'd20709;
          lut[4198] <= 16'd20755;
          lut[4199] <= 16'd20801;
          lut[4200] <= 16'd20845;
          lut[4201] <= 16'd20889;
          lut[4202] <= 16'd20932;
          lut[4203] <= 16'd20975;
          lut[4204] <= 16'd21016;
          lut[4205] <= 16'd21057;
          lut[4206] <= 16'd21098;
          lut[4207] <= 16'd21137;
          lut[4208] <= 16'd21176;
          lut[4209] <= 16'd21215;
          lut[4210] <= 16'd21252;
          lut[4211] <= 16'd21289;
          lut[4212] <= 16'd21326;
          lut[4213] <= 16'd21362;
          lut[4214] <= 16'd21397;
          lut[4215] <= 16'd21432;
          lut[4216] <= 16'd21466;
          lut[4217] <= 16'd21500;
          lut[4218] <= 16'd21533;
          lut[4219] <= 16'd21566;
          lut[4220] <= 16'd21598;
          lut[4221] <= 16'd21630;
          lut[4222] <= 16'd21661;
          lut[4223] <= 16'd21692;
          lut[4224] <= 0;
          lut[4225] <= 16'd496;
          lut[4226] <= 16'd992;
          lut[4227] <= 16'd1485;
          lut[4228] <= 16'd1976;
          lut[4229] <= 16'd2464;
          lut[4230] <= 16'd2947;
          lut[4231] <= 16'd3425;
          lut[4232] <= 16'd3897;
          lut[4233] <= 16'd4362;
          lut[4234] <= 16'd4821;
          lut[4235] <= 16'd5272;
          lut[4236] <= 16'd5714;
          lut[4237] <= 16'd6148;
          lut[4238] <= 16'd6574;
          lut[4239] <= 16'd6990;
          lut[4240] <= 16'd7397;
          lut[4241] <= 16'd7794;
          lut[4242] <= 16'd8181;
          lut[4243] <= 16'd8559;
          lut[4244] <= 16'd8927;
          lut[4245] <= 16'd9285;
          lut[4246] <= 16'd9634;
          lut[4247] <= 16'd9973;
          lut[4248] <= 16'd10302;
          lut[4249] <= 16'd10622;
          lut[4250] <= 16'd10933;
          lut[4251] <= 16'd11235;
          lut[4252] <= 16'd11528;
          lut[4253] <= 16'd11812;
          lut[4254] <= 16'd12088;
          lut[4255] <= 16'd12356;
          lut[4256] <= 16'd12616;
          lut[4257] <= 16'd12868;
          lut[4258] <= 16'd13112;
          lut[4259] <= 16'd13350;
          lut[4260] <= 16'd13580;
          lut[4261] <= 16'd13803;
          lut[4262] <= 16'd14020;
          lut[4263] <= 16'd14230;
          lut[4264] <= 16'd14434;
          lut[4265] <= 16'd14632;
          lut[4266] <= 16'd14825;
          lut[4267] <= 16'd15011;
          lut[4268] <= 16'd15193;
          lut[4269] <= 16'd15369;
          lut[4270] <= 16'd15540;
          lut[4271] <= 16'd15706;
          lut[4272] <= 16'd15868;
          lut[4273] <= 16'd16025;
          lut[4274] <= 16'd16178;
          lut[4275] <= 16'd16327;
          lut[4276] <= 16'd16471;
          lut[4277] <= 16'd16612;
          lut[4278] <= 16'd16748;
          lut[4279] <= 16'd16882;
          lut[4280] <= 16'd17011;
          lut[4281] <= 16'd17138;
          lut[4282] <= 16'd17261;
          lut[4283] <= 16'd17381;
          lut[4284] <= 16'd17497;
          lut[4285] <= 16'd17611;
          lut[4286] <= 16'd17722;
          lut[4287] <= 16'd17830;
          lut[4288] <= 16'd17936;
          lut[4289] <= 16'd18039;
          lut[4290] <= 16'd18140;
          lut[4291] <= 16'd18238;
          lut[4292] <= 16'd18333;
          lut[4293] <= 16'd18427;
          lut[4294] <= 16'd18518;
          lut[4295] <= 16'd18608;
          lut[4296] <= 16'd18695;
          lut[4297] <= 16'd18780;
          lut[4298] <= 16'd18863;
          lut[4299] <= 16'd18945;
          lut[4300] <= 16'd19024;
          lut[4301] <= 16'd19102;
          lut[4302] <= 16'd19178;
          lut[4303] <= 16'd19253;
          lut[4304] <= 16'd19326;
          lut[4305] <= 16'd19397;
          lut[4306] <= 16'd19467;
          lut[4307] <= 16'd19536;
          lut[4308] <= 16'd19603;
          lut[4309] <= 16'd19669;
          lut[4310] <= 16'd19733;
          lut[4311] <= 16'd19796;
          lut[4312] <= 16'd19858;
          lut[4313] <= 16'd19918;
          lut[4314] <= 16'd19978;
          lut[4315] <= 16'd20036;
          lut[4316] <= 16'd20093;
          lut[4317] <= 16'd20149;
          lut[4318] <= 16'd20204;
          lut[4319] <= 16'd20258;
          lut[4320] <= 16'd20311;
          lut[4321] <= 16'd20363;
          lut[4322] <= 16'd20414;
          lut[4323] <= 16'd20464;
          lut[4324] <= 16'd20514;
          lut[4325] <= 16'd20562;
          lut[4326] <= 16'd20609;
          lut[4327] <= 16'd20656;
          lut[4328] <= 16'd20702;
          lut[4329] <= 16'd20747;
          lut[4330] <= 16'd20791;
          lut[4331] <= 16'd20835;
          lut[4332] <= 16'd20877;
          lut[4333] <= 16'd20919;
          lut[4334] <= 16'd20961;
          lut[4335] <= 16'd21001;
          lut[4336] <= 16'd21041;
          lut[4337] <= 16'd21081;
          lut[4338] <= 16'd21119;
          lut[4339] <= 16'd21157;
          lut[4340] <= 16'd21195;
          lut[4341] <= 16'd21232;
          lut[4342] <= 16'd21268;
          lut[4343] <= 16'd21304;
          lut[4344] <= 16'd21339;
          lut[4345] <= 16'd21374;
          lut[4346] <= 16'd21408;
          lut[4347] <= 16'd21441;
          lut[4348] <= 16'd21474;
          lut[4349] <= 16'd21507;
          lut[4350] <= 16'd21539;
          lut[4351] <= 16'd21571;
          lut[4352] <= 0;
          lut[4353] <= 16'd482;
          lut[4354] <= 16'd963;
          lut[4355] <= 16'd1442;
          lut[4356] <= 16'd1919;
          lut[4357] <= 16'd2392;
          lut[4358] <= 16'd2862;
          lut[4359] <= 16'd3327;
          lut[4360] <= 16'd3786;
          lut[4361] <= 16'd4240;
          lut[4362] <= 16'd4687;
          lut[4363] <= 16'd5127;
          lut[4364] <= 16'd5559;
          lut[4365] <= 16'd5983;
          lut[4366] <= 16'd6400;
          lut[4367] <= 16'd6807;
          lut[4368] <= 16'd7206;
          lut[4369] <= 16'd7596;
          lut[4370] <= 16'd7977;
          lut[4371] <= 16'd8349;
          lut[4372] <= 16'd8712;
          lut[4373] <= 16'd9065;
          lut[4374] <= 16'd9409;
          lut[4375] <= 16'd9745;
          lut[4376] <= 16'd10071;
          lut[4377] <= 16'd10388;
          lut[4378] <= 16'd10696;
          lut[4379] <= 16'd10996;
          lut[4380] <= 16'd11287;
          lut[4381] <= 16'd11570;
          lut[4382] <= 16'd11845;
          lut[4383] <= 16'd12112;
          lut[4384] <= 16'd12372;
          lut[4385] <= 16'd12623;
          lut[4386] <= 16'd12868;
          lut[4387] <= 16'd13105;
          lut[4388] <= 16'd13336;
          lut[4389] <= 16'd13560;
          lut[4390] <= 16'd13777;
          lut[4391] <= 16'd13988;
          lut[4392] <= 16'd14193;
          lut[4393] <= 16'd14393;
          lut[4394] <= 16'd14586;
          lut[4395] <= 16'd14774;
          lut[4396] <= 16'd14957;
          lut[4397] <= 16'd15135;
          lut[4398] <= 16'd15307;
          lut[4399] <= 16'd15475;
          lut[4400] <= 16'd15639;
          lut[4401] <= 16'd15797;
          lut[4402] <= 16'd15952;
          lut[4403] <= 16'd16102;
          lut[4404] <= 16'd16248;
          lut[4405] <= 16'd16391;
          lut[4406] <= 16'd16529;
          lut[4407] <= 16'd16664;
          lut[4408] <= 16'd16796;
          lut[4409] <= 16'd16924;
          lut[4410] <= 16'd17049;
          lut[4411] <= 16'd17171;
          lut[4412] <= 16'd17289;
          lut[4413] <= 16'd17405;
          lut[4414] <= 16'd17518;
          lut[4415] <= 16'd17628;
          lut[4416] <= 16'd17735;
          lut[4417] <= 16'd17840;
          lut[4418] <= 16'd17942;
          lut[4419] <= 16'd18042;
          lut[4420] <= 16'd18140;
          lut[4421] <= 16'd18235;
          lut[4422] <= 16'd18328;
          lut[4423] <= 16'd18419;
          lut[4424] <= 16'd18508;
          lut[4425] <= 16'd18595;
          lut[4426] <= 16'd18679;
          lut[4427] <= 16'd18763;
          lut[4428] <= 16'd18844;
          lut[4429] <= 16'd18923;
          lut[4430] <= 16'd19001;
          lut[4431] <= 16'd19077;
          lut[4432] <= 16'd19152;
          lut[4433] <= 16'd19225;
          lut[4434] <= 16'd19296;
          lut[4435] <= 16'd19366;
          lut[4436] <= 16'd19435;
          lut[4437] <= 16'd19502;
          lut[4438] <= 16'd19568;
          lut[4439] <= 16'd19632;
          lut[4440] <= 16'd19695;
          lut[4441] <= 16'd19757;
          lut[4442] <= 16'd19818;
          lut[4443] <= 16'd19878;
          lut[4444] <= 16'd19936;
          lut[4445] <= 16'd19993;
          lut[4446] <= 16'd20050;
          lut[4447] <= 16'd20105;
          lut[4448] <= 16'd20159;
          lut[4449] <= 16'd20212;
          lut[4450] <= 16'd20265;
          lut[4451] <= 16'd20316;
          lut[4452] <= 16'd20366;
          lut[4453] <= 16'd20416;
          lut[4454] <= 16'd20464;
          lut[4455] <= 16'd20512;
          lut[4456] <= 16'd20559;
          lut[4457] <= 16'd20605;
          lut[4458] <= 16'd20651;
          lut[4459] <= 16'd20695;
          lut[4460] <= 16'd20739;
          lut[4461] <= 16'd20782;
          lut[4462] <= 16'd20824;
          lut[4463] <= 16'd20866;
          lut[4464] <= 16'd20907;
          lut[4465] <= 16'd20947;
          lut[4466] <= 16'd20987;
          lut[4467] <= 16'd21026;
          lut[4468] <= 16'd21065;
          lut[4469] <= 16'd21102;
          lut[4470] <= 16'd21140;
          lut[4471] <= 16'd21176;
          lut[4472] <= 16'd21212;
          lut[4473] <= 16'd21248;
          lut[4474] <= 16'd21283;
          lut[4475] <= 16'd21317;
          lut[4476] <= 16'd21351;
          lut[4477] <= 16'd21385;
          lut[4478] <= 16'd21418;
          lut[4479] <= 16'd21450;
          lut[4480] <= 0;
          lut[4481] <= 16'd468;
          lut[4482] <= 16'd935;
          lut[4483] <= 16'd1401;
          lut[4484] <= 16'd1864;
          lut[4485] <= 16'd2325;
          lut[4486] <= 16'd2782;
          lut[4487] <= 16'd3234;
          lut[4488] <= 16'd3682;
          lut[4489] <= 16'd4124;
          lut[4490] <= 16'd4560;
          lut[4491] <= 16'd4989;
          lut[4492] <= 16'd5412;
          lut[4493] <= 16'd5827;
          lut[4494] <= 16'd6234;
          lut[4495] <= 16'd6634;
          lut[4496] <= 16'd7025;
          lut[4497] <= 16'd7408;
          lut[4498] <= 16'd7783;
          lut[4499] <= 16'd8148;
          lut[4500] <= 16'd8506;
          lut[4501] <= 16'd8854;
          lut[4502] <= 16'd9194;
          lut[4503] <= 16'd9525;
          lut[4504] <= 16'd9848;
          lut[4505] <= 16'd10162;
          lut[4506] <= 16'd10468;
          lut[4507] <= 16'd10766;
          lut[4508] <= 16'd11055;
          lut[4509] <= 16'd11336;
          lut[4510] <= 16'd11610;
          lut[4511] <= 16'd11876;
          lut[4512] <= 16'd12135;
          lut[4513] <= 16'd12386;
          lut[4514] <= 16'd12631;
          lut[4515] <= 16'd12868;
          lut[4516] <= 16'd13099;
          lut[4517] <= 16'd13323;
          lut[4518] <= 16'd13541;
          lut[4519] <= 16'd13753;
          lut[4520] <= 16'd13959;
          lut[4521] <= 16'd14159;
          lut[4522] <= 16'd14353;
          lut[4523] <= 16'd14543;
          lut[4524] <= 16'd14726;
          lut[4525] <= 16'd14905;
          lut[4526] <= 16'd15079;
          lut[4527] <= 16'd15249;
          lut[4528] <= 16'd15413;
          lut[4529] <= 16'd15574;
          lut[4530] <= 16'd15730;
          lut[4531] <= 16'd15882;
          lut[4532] <= 16'd16030;
          lut[4533] <= 16'd16174;
          lut[4534] <= 16'd16314;
          lut[4535] <= 16'd16451;
          lut[4536] <= 16'd16584;
          lut[4537] <= 16'd16714;
          lut[4538] <= 16'd16840;
          lut[4539] <= 16'd16964;
          lut[4540] <= 16'd17084;
          lut[4541] <= 16'd17201;
          lut[4542] <= 16'd17316;
          lut[4543] <= 16'd17428;
          lut[4544] <= 16'd17537;
          lut[4545] <= 16'd17643;
          lut[4546] <= 16'd17747;
          lut[4547] <= 16'd17849;
          lut[4548] <= 16'd17948;
          lut[4549] <= 16'd18045;
          lut[4550] <= 16'd18140;
          lut[4551] <= 16'd18232;
          lut[4552] <= 16'd18323;
          lut[4553] <= 16'd18411;
          lut[4554] <= 16'd18498;
          lut[4555] <= 16'd18582;
          lut[4556] <= 16'd18665;
          lut[4557] <= 16'd18746;
          lut[4558] <= 16'd18825;
          lut[4559] <= 16'd18903;
          lut[4560] <= 16'd18979;
          lut[4561] <= 16'd19053;
          lut[4562] <= 16'd19126;
          lut[4563] <= 16'd19198;
          lut[4564] <= 16'd19268;
          lut[4565] <= 16'd19336;
          lut[4566] <= 16'd19403;
          lut[4567] <= 16'd19469;
          lut[4568] <= 16'd19534;
          lut[4569] <= 16'd19597;
          lut[4570] <= 16'd19659;
          lut[4571] <= 16'd19720;
          lut[4572] <= 16'd19780;
          lut[4573] <= 16'd19839;
          lut[4574] <= 16'd19896;
          lut[4575] <= 16'd19953;
          lut[4576] <= 16'd20008;
          lut[4577] <= 16'd20062;
          lut[4578] <= 16'd20116;
          lut[4579] <= 16'd20168;
          lut[4580] <= 16'd20220;
          lut[4581] <= 16'd20270;
          lut[4582] <= 16'd20320;
          lut[4583] <= 16'd20369;
          lut[4584] <= 16'd20417;
          lut[4585] <= 16'd20464;
          lut[4586] <= 16'd20511;
          lut[4587] <= 16'd20556;
          lut[4588] <= 16'd20601;
          lut[4589] <= 16'd20645;
          lut[4590] <= 16'd20689;
          lut[4591] <= 16'd20731;
          lut[4592] <= 16'd20773;
          lut[4593] <= 16'd20815;
          lut[4594] <= 16'd20855;
          lut[4595] <= 16'd20895;
          lut[4596] <= 16'd20935;
          lut[4597] <= 16'd20974;
          lut[4598] <= 16'd21012;
          lut[4599] <= 16'd21049;
          lut[4600] <= 16'd21086;
          lut[4601] <= 16'd21123;
          lut[4602] <= 16'd21159;
          lut[4603] <= 16'd21194;
          lut[4604] <= 16'd21229;
          lut[4605] <= 16'd21263;
          lut[4606] <= 16'd21297;
          lut[4607] <= 16'd21330;
          lut[4608] <= 0;
          lut[4609] <= 16'd455;
          lut[4610] <= 16'd909;
          lut[4611] <= 16'd1362;
          lut[4612] <= 16'd1813;
          lut[4613] <= 16'd2261;
          lut[4614] <= 16'd2706;
          lut[4615] <= 16'd3147;
          lut[4616] <= 16'd3583;
          lut[4617] <= 16'd4014;
          lut[4618] <= 16'd4439;
          lut[4619] <= 16'd4859;
          lut[4620] <= 16'd5272;
          lut[4621] <= 16'd5678;
          lut[4622] <= 16'd6077;
          lut[4623] <= 16'd6468;
          lut[4624] <= 16'd6852;
          lut[4625] <= 16'd7228;
          lut[4626] <= 16'd7596;
          lut[4627] <= 16'd7956;
          lut[4628] <= 16'd8308;
          lut[4629] <= 16'd8652;
          lut[4630] <= 16'd8987;
          lut[4631] <= 16'd9315;
          lut[4632] <= 16'd9634;
          lut[4633] <= 16'd9945;
          lut[4634] <= 16'd10248;
          lut[4635] <= 16'd10543;
          lut[4636] <= 16'd10831;
          lut[4637] <= 16'd11110;
          lut[4638] <= 16'd11383;
          lut[4639] <= 16'd11648;
          lut[4640] <= 16'd11905;
          lut[4641] <= 16'd12156;
          lut[4642] <= 16'd12400;
          lut[4643] <= 16'd12637;
          lut[4644] <= 16'd12868;
          lut[4645] <= 16'd13092;
          lut[4646] <= 16'd13311;
          lut[4647] <= 16'd13523;
          lut[4648] <= 16'd13729;
          lut[4649] <= 16'd13930;
          lut[4650] <= 16'd14126;
          lut[4651] <= 16'd14316;
          lut[4652] <= 16'd14501;
          lut[4653] <= 16'd14681;
          lut[4654] <= 16'd14856;
          lut[4655] <= 16'd15027;
          lut[4656] <= 16'd15193;
          lut[4657] <= 16'd15354;
          lut[4658] <= 16'd15512;
          lut[4659] <= 16'd15665;
          lut[4660] <= 16'd15815;
          lut[4661] <= 16'd15960;
          lut[4662] <= 16'd16102;
          lut[4663] <= 16'd16240;
          lut[4664] <= 16'd16375;
          lut[4665] <= 16'd16507;
          lut[4666] <= 16'd16635;
          lut[4667] <= 16'd16760;
          lut[4668] <= 16'd16882;
          lut[4669] <= 16'd17001;
          lut[4670] <= 16'd17117;
          lut[4671] <= 16'd17230;
          lut[4672] <= 16'd17341;
          lut[4673] <= 16'd17449;
          lut[4674] <= 16'd17555;
          lut[4675] <= 16'd17658;
          lut[4676] <= 16'd17759;
          lut[4677] <= 16'd17857;
          lut[4678] <= 16'd17953;
          lut[4679] <= 16'd18047;
          lut[4680] <= 16'd18140;
          lut[4681] <= 16'd18230;
          lut[4682] <= 16'd18318;
          lut[4683] <= 16'd18404;
          lut[4684] <= 16'd18488;
          lut[4685] <= 16'd18571;
          lut[4686] <= 16'd18651;
          lut[4687] <= 16'd18730;
          lut[4688] <= 16'd18808;
          lut[4689] <= 16'd18884;
          lut[4690] <= 16'd18958;
          lut[4691] <= 16'd19031;
          lut[4692] <= 16'd19102;
          lut[4693] <= 16'd19172;
          lut[4694] <= 16'd19241;
          lut[4695] <= 16'd19308;
          lut[4696] <= 16'd19374;
          lut[4697] <= 16'd19438;
          lut[4698] <= 16'd19502;
          lut[4699] <= 16'd19564;
          lut[4700] <= 16'd19625;
          lut[4701] <= 16'd19685;
          lut[4702] <= 16'd19744;
          lut[4703] <= 16'd19801;
          lut[4704] <= 16'd19858;
          lut[4705] <= 16'd19913;
          lut[4706] <= 16'd19968;
          lut[4707] <= 16'd20022;
          lut[4708] <= 16'd20074;
          lut[4709] <= 16'd20126;
          lut[4710] <= 16'd20177;
          lut[4711] <= 16'd20227;
          lut[4712] <= 16'd20276;
          lut[4713] <= 16'd20324;
          lut[4714] <= 16'd20372;
          lut[4715] <= 16'd20418;
          lut[4716] <= 16'd20464;
          lut[4717] <= 16'd20510;
          lut[4718] <= 16'd20554;
          lut[4719] <= 16'd20598;
          lut[4720] <= 16'd20641;
          lut[4721] <= 16'd20683;
          lut[4722] <= 16'd20724;
          lut[4723] <= 16'd20765;
          lut[4724] <= 16'd20806;
          lut[4725] <= 16'd20845;
          lut[4726] <= 16'd20884;
          lut[4727] <= 16'd20923;
          lut[4728] <= 16'd20961;
          lut[4729] <= 16'd20998;
          lut[4730] <= 16'd21035;
          lut[4731] <= 16'd21071;
          lut[4732] <= 16'd21107;
          lut[4733] <= 16'd21142;
          lut[4734] <= 16'd21176;
          lut[4735] <= 16'd21210;
          lut[4736] <= 0;
          lut[4737] <= 16'd443;
          lut[4738] <= 16'd885;
          lut[4739] <= 16'd1326;
          lut[4740] <= 16'd1764;
          lut[4741] <= 16'd2201;
          lut[4742] <= 16'd2634;
          lut[4743] <= 16'd3063;
          lut[4744] <= 16'd3489;
          lut[4745] <= 16'd3909;
          lut[4746] <= 16'd4325;
          lut[4747] <= 16'd4735;
          lut[4748] <= 16'd5138;
          lut[4749] <= 16'd5536;
          lut[4750] <= 16'd5927;
          lut[4751] <= 16'd6310;
          lut[4752] <= 16'd6687;
          lut[4753] <= 16'd7056;
          lut[4754] <= 16'd7418;
          lut[4755] <= 16'd7773;
          lut[4756] <= 16'd8119;
          lut[4757] <= 16'd8458;
          lut[4758] <= 16'd8789;
          lut[4759] <= 16'd9112;
          lut[4760] <= 16'd9428;
          lut[4761] <= 16'd9736;
          lut[4762] <= 16'd10036;
          lut[4763] <= 16'd10328;
          lut[4764] <= 16'd10614;
          lut[4765] <= 16'd10892;
          lut[4766] <= 16'd11162;
          lut[4767] <= 16'd11426;
          lut[4768] <= 16'd11683;
          lut[4769] <= 16'd11933;
          lut[4770] <= 16'd12176;
          lut[4771] <= 16'd12413;
          lut[4772] <= 16'd12644;
          lut[4773] <= 16'd12868;
          lut[4774] <= 16'd13086;
          lut[4775] <= 16'd13299;
          lut[4776] <= 16'd13506;
          lut[4777] <= 16'd13707;
          lut[4778] <= 16'd13904;
          lut[4779] <= 16'd14094;
          lut[4780] <= 16'd14280;
          lut[4781] <= 16'd14461;
          lut[4782] <= 16'd14638;
          lut[4783] <= 16'd14809;
          lut[4784] <= 16'd14977;
          lut[4785] <= 16'd15139;
          lut[4786] <= 16'd15298;
          lut[4787] <= 16'd15453;
          lut[4788] <= 16'd15604;
          lut[4789] <= 16'd15751;
          lut[4790] <= 16'd15894;
          lut[4791] <= 16'd16034;
          lut[4792] <= 16'd16170;
          lut[4793] <= 16'd16303;
          lut[4794] <= 16'd16432;
          lut[4795] <= 16'd16559;
          lut[4796] <= 16'd16682;
          lut[4797] <= 16'd16803;
          lut[4798] <= 16'd16921;
          lut[4799] <= 16'd17036;
          lut[4800] <= 16'd17148;
          lut[4801] <= 16'd17257;
          lut[4802] <= 16'd17365;
          lut[4803] <= 16'd17469;
          lut[4804] <= 16'd17572;
          lut[4805] <= 16'd17672;
          lut[4806] <= 16'd17769;
          lut[4807] <= 16'd17865;
          lut[4808] <= 16'd17958;
          lut[4809] <= 16'd18050;
          lut[4810] <= 16'd18140;
          lut[4811] <= 16'd18227;
          lut[4812] <= 16'd18313;
          lut[4813] <= 16'd18397;
          lut[4814] <= 16'd18479;
          lut[4815] <= 16'd18560;
          lut[4816] <= 16'd18638;
          lut[4817] <= 16'd18716;
          lut[4818] <= 16'd18791;
          lut[4819] <= 16'd18865;
          lut[4820] <= 16'd18938;
          lut[4821] <= 16'd19009;
          lut[4822] <= 16'd19079;
          lut[4823] <= 16'd19148;
          lut[4824] <= 16'd19215;
          lut[4825] <= 16'd19281;
          lut[4826] <= 16'd19345;
          lut[4827] <= 16'd19409;
          lut[4828] <= 16'd19471;
          lut[4829] <= 16'd19532;
          lut[4830] <= 16'd19592;
          lut[4831] <= 16'd19651;
          lut[4832] <= 16'd19709;
          lut[4833] <= 16'd19765;
          lut[4834] <= 16'd19821;
          lut[4835] <= 16'd19876;
          lut[4836] <= 16'd19930;
          lut[4837] <= 16'd19983;
          lut[4838] <= 16'd20035;
          lut[4839] <= 16'd20086;
          lut[4840] <= 16'd20136;
          lut[4841] <= 16'd20185;
          lut[4842] <= 16'd20234;
          lut[4843] <= 16'd20281;
          lut[4844] <= 16'd20328;
          lut[4845] <= 16'd20374;
          lut[4846] <= 16'd20420;
          lut[4847] <= 16'd20464;
          lut[4848] <= 16'd20508;
          lut[4849] <= 16'd20552;
          lut[4850] <= 16'd20594;
          lut[4851] <= 16'd20636;
          lut[4852] <= 16'd20677;
          lut[4853] <= 16'd20718;
          lut[4854] <= 16'd20758;
          lut[4855] <= 16'd20797;
          lut[4856] <= 16'd20836;
          lut[4857] <= 16'd20874;
          lut[4858] <= 16'd20911;
          lut[4859] <= 16'd20948;
          lut[4860] <= 16'd20985;
          lut[4861] <= 16'd21021;
          lut[4862] <= 16'd21056;
          lut[4863] <= 16'd21091;
          lut[4864] <= 0;
          lut[4865] <= 16'd431;
          lut[4866] <= 16'd862;
          lut[4867] <= 16'd1291;
          lut[4868] <= 16'd1718;
          lut[4869] <= 16'd2143;
          lut[4870] <= 16'd2566;
          lut[4871] <= 16'd2985;
          lut[4872] <= 16'd3400;
          lut[4873] <= 16'd3810;
          lut[4874] <= 16'd4216;
          lut[4875] <= 16'd4617;
          lut[4876] <= 16'd5012;
          lut[4877] <= 16'd5401;
          lut[4878] <= 16'd5783;
          lut[4879] <= 16'd6160;
          lut[4880] <= 16'd6529;
          lut[4881] <= 16'd6892;
          lut[4882] <= 16'd7248;
          lut[4883] <= 16'd7596;
          lut[4884] <= 16'd7938;
          lut[4885] <= 16'd8272;
          lut[4886] <= 16'd8598;
          lut[4887] <= 16'd8917;
          lut[4888] <= 16'd9229;
          lut[4889] <= 16'd9534;
          lut[4890] <= 16'd9831;
          lut[4891] <= 16'd10121;
          lut[4892] <= 16'd10404;
          lut[4893] <= 16'd10680;
          lut[4894] <= 16'd10949;
          lut[4895] <= 16'd11211;
          lut[4896] <= 16'd11467;
          lut[4897] <= 16'd11716;
          lut[4898] <= 16'd11959;
          lut[4899] <= 16'd12195;
          lut[4900] <= 16'd12425;
          lut[4901] <= 16'd12650;
          lut[4902] <= 16'd12868;
          lut[4903] <= 16'd13081;
          lut[4904] <= 16'd13288;
          lut[4905] <= 16'd13490;
          lut[4906] <= 16'd13686;
          lut[4907] <= 16'd13878;
          lut[4908] <= 16'd14065;
          lut[4909] <= 16'd14246;
          lut[4910] <= 16'd14424;
          lut[4911] <= 16'd14596;
          lut[4912] <= 16'd14765;
          lut[4913] <= 16'd14929;
          lut[4914] <= 16'd15088;
          lut[4915] <= 16'd15244;
          lut[4916] <= 16'd15396;
          lut[4917] <= 16'd15545;
          lut[4918] <= 16'd15689;
          lut[4919] <= 16'd15830;
          lut[4920] <= 16'd15968;
          lut[4921] <= 16'd16102;
          lut[4922] <= 16'd16233;
          lut[4923] <= 16'd16361;
          lut[4924] <= 16'd16486;
          lut[4925] <= 16'd16608;
          lut[4926] <= 16'd16727;
          lut[4927] <= 16'd16844;
          lut[4928] <= 16'd16957;
          lut[4929] <= 16'd17068;
          lut[4930] <= 16'd17177;
          lut[4931] <= 16'd17283;
          lut[4932] <= 16'd17387;
          lut[4933] <= 16'd17488;
          lut[4934] <= 16'd17587;
          lut[4935] <= 16'd17685;
          lut[4936] <= 16'd17779;
          lut[4937] <= 16'd17872;
          lut[4938] <= 16'd17963;
          lut[4939] <= 16'd18052;
          lut[4940] <= 16'd18140;
          lut[4941] <= 16'd18225;
          lut[4942] <= 16'd18308;
          lut[4943] <= 16'd18390;
          lut[4944] <= 16'd18470;
          lut[4945] <= 16'd18549;
          lut[4946] <= 16'd18626;
          lut[4947] <= 16'd18702;
          lut[4948] <= 16'd18775;
          lut[4949] <= 16'd18848;
          lut[4950] <= 16'd18919;
          lut[4951] <= 16'd18989;
          lut[4952] <= 16'd19057;
          lut[4953] <= 16'd19124;
          lut[4954] <= 16'd19190;
          lut[4955] <= 16'd19255;
          lut[4956] <= 16'd19318;
          lut[4957] <= 16'd19381;
          lut[4958] <= 16'd19442;
          lut[4959] <= 16'd19502;
          lut[4960] <= 16'd19561;
          lut[4961] <= 16'd19619;
          lut[4962] <= 16'd19675;
          lut[4963] <= 16'd19731;
          lut[4964] <= 16'd19786;
          lut[4965] <= 16'd19840;
          lut[4966] <= 16'd19893;
          lut[4967] <= 16'd19945;
          lut[4968] <= 16'd19996;
          lut[4969] <= 16'd20047;
          lut[4970] <= 16'd20096;
          lut[4971] <= 16'd20145;
          lut[4972] <= 16'd20193;
          lut[4973] <= 16'd20240;
          lut[4974] <= 16'd20286;
          lut[4975] <= 16'd20332;
          lut[4976] <= 16'd20377;
          lut[4977] <= 16'd20421;
          lut[4978] <= 16'd20464;
          lut[4979] <= 16'd20507;
          lut[4980] <= 16'd20549;
          lut[4981] <= 16'd20591;
          lut[4982] <= 16'd20632;
          lut[4983] <= 16'd20672;
          lut[4984] <= 16'd20711;
          lut[4985] <= 16'd20750;
          lut[4986] <= 16'd20789;
          lut[4987] <= 16'd20827;
          lut[4988] <= 16'd20864;
          lut[4989] <= 16'd20901;
          lut[4990] <= 16'd20937;
          lut[4991] <= 16'd20973;
          lut[4992] <= 0;
          lut[4993] <= 16'd420;
          lut[4994] <= 16'd839;
          lut[4995] <= 16'd1258;
          lut[4996] <= 16'd1675;
          lut[4997] <= 16'd2089;
          lut[4998] <= 16'd2501;
          lut[4999] <= 16'd2910;
          lut[5000] <= 16'd3315;
          lut[5001] <= 16'd3716;
          lut[5002] <= 16'd4112;
          lut[5003] <= 16'd4504;
          lut[5004] <= 16'd4891;
          lut[5005] <= 16'd5272;
          lut[5006] <= 16'd5647;
          lut[5007] <= 16'd6016;
          lut[5008] <= 16'd6379;
          lut[5009] <= 16'd6735;
          lut[5010] <= 16'd7085;
          lut[5011] <= 16'd7428;
          lut[5012] <= 16'd7764;
          lut[5013] <= 16'd8093;
          lut[5014] <= 16'd8415;
          lut[5015] <= 16'd8730;
          lut[5016] <= 16'd9038;
          lut[5017] <= 16'd9340;
          lut[5018] <= 16'd9634;
          lut[5019] <= 16'd9921;
          lut[5020] <= 16'd10202;
          lut[5021] <= 16'd10476;
          lut[5022] <= 16'd10743;
          lut[5023] <= 16'd11004;
          lut[5024] <= 16'd11258;
          lut[5025] <= 16'd11506;
          lut[5026] <= 16'd11748;
          lut[5027] <= 16'd11983;
          lut[5028] <= 16'd12213;
          lut[5029] <= 16'd12437;
          lut[5030] <= 16'd12655;
          lut[5031] <= 16'd12868;
          lut[5032] <= 16'd13075;
          lut[5033] <= 16'd13277;
          lut[5034] <= 16'd13475;
          lut[5035] <= 16'd13667;
          lut[5036] <= 16'd13854;
          lut[5037] <= 16'd14036;
          lut[5038] <= 16'd14214;
          lut[5039] <= 16'd14388;
          lut[5040] <= 16'd14557;
          lut[5041] <= 16'd14722;
          lut[5042] <= 16'd14883;
          lut[5043] <= 16'd15040;
          lut[5044] <= 16'd15193;
          lut[5045] <= 16'd15342;
          lut[5046] <= 16'd15488;
          lut[5047] <= 16'd15630;
          lut[5048] <= 16'd15769;
          lut[5049] <= 16'd15905;
          lut[5050] <= 16'd16037;
          lut[5051] <= 16'd16166;
          lut[5052] <= 16'd16293;
          lut[5053] <= 16'd16416;
          lut[5054] <= 16'd16536;
          lut[5055] <= 16'd16654;
          lut[5056] <= 16'd16769;
          lut[5057] <= 16'd16882;
          lut[5058] <= 16'd16992;
          lut[5059] <= 16'd17099;
          lut[5060] <= 16'd17204;
          lut[5061] <= 16'd17307;
          lut[5062] <= 16'd17408;
          lut[5063] <= 16'd17506;
          lut[5064] <= 16'd17603;
          lut[5065] <= 16'd17697;
          lut[5066] <= 16'd17789;
          lut[5067] <= 16'd17879;
          lut[5068] <= 16'd17968;
          lut[5069] <= 16'd18055;
          lut[5070] <= 16'd18140;
          lut[5071] <= 16'd18223;
          lut[5072] <= 16'd18304;
          lut[5073] <= 16'd18384;
          lut[5074] <= 16'd18462;
          lut[5075] <= 16'd18539;
          lut[5076] <= 16'd18614;
          lut[5077] <= 16'd18688;
          lut[5078] <= 16'd18760;
          lut[5079] <= 16'd18831;
          lut[5080] <= 16'd18901;
          lut[5081] <= 16'd18969;
          lut[5082] <= 16'd19036;
          lut[5083] <= 16'd19102;
          lut[5084] <= 16'd19167;
          lut[5085] <= 16'd19230;
          lut[5086] <= 16'd19292;
          lut[5087] <= 16'd19354;
          lut[5088] <= 16'd19414;
          lut[5089] <= 16'd19473;
          lut[5090] <= 16'd19531;
          lut[5091] <= 16'd19587;
          lut[5092] <= 16'd19643;
          lut[5093] <= 16'd19698;
          lut[5094] <= 16'd19752;
          lut[5095] <= 16'd19806;
          lut[5096] <= 16'd19858;
          lut[5097] <= 16'd19909;
          lut[5098] <= 16'd19960;
          lut[5099] <= 16'd20009;
          lut[5100] <= 16'd20058;
          lut[5101] <= 16'd20106;
          lut[5102] <= 16'd20154;
          lut[5103] <= 16'd20200;
          lut[5104] <= 16'd20246;
          lut[5105] <= 16'd20291;
          lut[5106] <= 16'd20335;
          lut[5107] <= 16'd20379;
          lut[5108] <= 16'd20422;
          lut[5109] <= 16'd20464;
          lut[5110] <= 16'd20506;
          lut[5111] <= 16'd20547;
          lut[5112] <= 16'd20588;
          lut[5113] <= 16'd20627;
          lut[5114] <= 16'd20667;
          lut[5115] <= 16'd20705;
          lut[5116] <= 16'd20743;
          lut[5117] <= 16'd20781;
          lut[5118] <= 16'd20818;
          lut[5119] <= 16'd20854;
          lut[5120] <= 0;
          lut[5121] <= 16'd410;
          lut[5122] <= 16'd819;
          lut[5123] <= 16'd1227;
          lut[5124] <= 16'd1633;
          lut[5125] <= 16'd2037;
          lut[5126] <= 16'd2439;
          lut[5127] <= 16'd2838;
          lut[5128] <= 16'd3234;
          lut[5129] <= 16'd3626;
          lut[5130] <= 16'd4014;
          lut[5131] <= 16'd4397;
          lut[5132] <= 16'd4775;
          lut[5133] <= 16'd5148;
          lut[5134] <= 16'd5516;
          lut[5135] <= 16'd5878;
          lut[5136] <= 16'd6234;
          lut[5137] <= 16'd6584;
          lut[5138] <= 16'd6928;
          lut[5139] <= 16'd7265;
          lut[5140] <= 16'd7596;
          lut[5141] <= 16'd7921;
          lut[5142] <= 16'd8239;
          lut[5143] <= 16'd8550;
          lut[5144] <= 16'd8854;
          lut[5145] <= 16'd9152;
          lut[5146] <= 16'd9443;
          lut[5147] <= 16'd9728;
          lut[5148] <= 16'd10006;
          lut[5149] <= 16'd10278;
          lut[5150] <= 16'd10543;
          lut[5151] <= 16'd10802;
          lut[5152] <= 16'd11055;
          lut[5153] <= 16'd11302;
          lut[5154] <= 16'd11542;
          lut[5155] <= 16'd11777;
          lut[5156] <= 16'd12006;
          lut[5157] <= 16'd12230;
          lut[5158] <= 16'd12448;
          lut[5159] <= 16'd12661;
          lut[5160] <= 16'd12868;
          lut[5161] <= 16'd13070;
          lut[5162] <= 16'd13267;
          lut[5163] <= 16'd13460;
          lut[5164] <= 16'd13648;
          lut[5165] <= 16'd13831;
          lut[5166] <= 16'd14009;
          lut[5167] <= 16'd14183;
          lut[5168] <= 16'd14353;
          lut[5169] <= 16'd14519;
          lut[5170] <= 16'd14681;
          lut[5171] <= 16'd14839;
          lut[5172] <= 16'd14993;
          lut[5173] <= 16'd15143;
          lut[5174] <= 16'd15290;
          lut[5175] <= 16'd15434;
          lut[5176] <= 16'd15574;
          lut[5177] <= 16'd15711;
          lut[5178] <= 16'd15844;
          lut[5179] <= 16'd15975;
          lut[5180] <= 16'd16102;
          lut[5181] <= 16'd16227;
          lut[5182] <= 16'd16348;
          lut[5183] <= 16'd16467;
          lut[5184] <= 16'd16584;
          lut[5185] <= 16'd16698;
          lut[5186] <= 16'd16809;
          lut[5187] <= 16'd16918;
          lut[5188] <= 16'd17024;
          lut[5189] <= 16'd17128;
          lut[5190] <= 16'd17230;
          lut[5191] <= 16'd17330;
          lut[5192] <= 16'd17428;
          lut[5193] <= 16'd17523;
          lut[5194] <= 16'd17617;
          lut[5195] <= 16'd17708;
          lut[5196] <= 16'd17798;
          lut[5197] <= 16'd17886;
          lut[5198] <= 16'd17972;
          lut[5199] <= 16'd18057;
          lut[5200] <= 16'd18140;
          lut[5201] <= 16'd18221;
          lut[5202] <= 16'd18300;
          lut[5203] <= 16'd18378;
          lut[5204] <= 16'd18455;
          lut[5205] <= 16'd18530;
          lut[5206] <= 16'd18603;
          lut[5207] <= 16'd18675;
          lut[5208] <= 16'd18746;
          lut[5209] <= 16'd18816;
          lut[5210] <= 16'd18884;
          lut[5211] <= 16'd18951;
          lut[5212] <= 16'd19016;
          lut[5213] <= 16'd19081;
          lut[5214] <= 16'd19144;
          lut[5215] <= 16'd19207;
          lut[5216] <= 16'd19268;
          lut[5217] <= 16'd19328;
          lut[5218] <= 16'd19387;
          lut[5219] <= 16'd19445;
          lut[5220] <= 16'd19502;
          lut[5221] <= 16'd19558;
          lut[5222] <= 16'd19613;
          lut[5223] <= 16'd19667;
          lut[5224] <= 16'd19720;
          lut[5225] <= 16'd19772;
          lut[5226] <= 16'd19824;
          lut[5227] <= 16'd19875;
          lut[5228] <= 16'd19924;
          lut[5229] <= 16'd19973;
          lut[5230] <= 16'd20022;
          lut[5231] <= 16'd20069;
          lut[5232] <= 16'd20116;
          lut[5233] <= 16'd20162;
          lut[5234] <= 16'd20207;
          lut[5235] <= 16'd20252;
          lut[5236] <= 16'd20295;
          lut[5237] <= 16'd20339;
          lut[5238] <= 16'd20381;
          lut[5239] <= 16'd20423;
          lut[5240] <= 16'd20464;
          lut[5241] <= 16'd20505;
          lut[5242] <= 16'd20545;
          lut[5243] <= 16'd20585;
          lut[5244] <= 16'd20623;
          lut[5245] <= 16'd20662;
          lut[5246] <= 16'd20700;
          lut[5247] <= 16'd20737;
          lut[5248] <= 0;
          lut[5249] <= 16'd400;
          lut[5250] <= 16'd799;
          lut[5251] <= 16'd1197;
          lut[5252] <= 16'd1593;
          lut[5253] <= 16'd1988;
          lut[5254] <= 16'd2381;
          lut[5255] <= 16'd2771;
          lut[5256] <= 16'd3157;
          lut[5257] <= 16'd3540;
          lut[5258] <= 16'd3920;
          lut[5259] <= 16'd4295;
          lut[5260] <= 16'd4665;
          lut[5261] <= 16'd5031;
          lut[5262] <= 16'd5391;
          lut[5263] <= 16'd5746;
          lut[5264] <= 16'd6096;
          lut[5265] <= 16'd6440;
          lut[5266] <= 16'd6778;
          lut[5267] <= 16'd7110;
          lut[5268] <= 16'd7436;
          lut[5269] <= 16'd7755;
          lut[5270] <= 16'd8069;
          lut[5271] <= 16'd8376;
          lut[5272] <= 16'd8677;
          lut[5273] <= 16'd8971;
          lut[5274] <= 16'd9259;
          lut[5275] <= 16'd9541;
          lut[5276] <= 16'd9817;
          lut[5277] <= 16'd10086;
          lut[5278] <= 16'd10350;
          lut[5279] <= 16'd10607;
          lut[5280] <= 16'd10858;
          lut[5281] <= 16'd11104;
          lut[5282] <= 16'd11343;
          lut[5283] <= 16'd11577;
          lut[5284] <= 16'd11806;
          lut[5285] <= 16'd12028;
          lut[5286] <= 16'd12246;
          lut[5287] <= 16'd12458;
          lut[5288] <= 16'd12666;
          lut[5289] <= 16'd12868;
          lut[5290] <= 16'd13065;
          lut[5291] <= 16'd13258;
          lut[5292] <= 16'd13446;
          lut[5293] <= 16'd13629;
          lut[5294] <= 16'd13809;
          lut[5295] <= 16'd13983;
          lut[5296] <= 16'd14154;
          lut[5297] <= 16'd14321;
          lut[5298] <= 16'd14483;
          lut[5299] <= 16'd14642;
          lut[5300] <= 16'd14797;
          lut[5301] <= 16'd14948;
          lut[5302] <= 16'd15096;
          lut[5303] <= 16'd15241;
          lut[5304] <= 16'd15382;
          lut[5305] <= 16'd15520;
          lut[5306] <= 16'd15654;
          lut[5307] <= 16'd15786;
          lut[5308] <= 16'd15914;
          lut[5309] <= 16'd16040;
          lut[5310] <= 16'd16163;
          lut[5311] <= 16'd16283;
          lut[5312] <= 16'd16401;
          lut[5313] <= 16'd16516;
          lut[5314] <= 16'd16629;
          lut[5315] <= 16'd16739;
          lut[5316] <= 16'd16846;
          lut[5317] <= 16'd16952;
          lut[5318] <= 16'd17055;
          lut[5319] <= 16'd17156;
          lut[5320] <= 16'd17255;
          lut[5321] <= 16'd17352;
          lut[5322] <= 16'd17446;
          lut[5323] <= 16'd17539;
          lut[5324] <= 16'd17630;
          lut[5325] <= 16'd17720;
          lut[5326] <= 16'd17807;
          lut[5327] <= 16'd17893;
          lut[5328] <= 16'd17977;
          lut[5329] <= 16'd18059;
          lut[5330] <= 16'd18140;
          lut[5331] <= 16'd18219;
          lut[5332] <= 16'd18296;
          lut[5333] <= 16'd18372;
          lut[5334] <= 16'd18447;
          lut[5335] <= 16'd18520;
          lut[5336] <= 16'd18592;
          lut[5337] <= 16'd18663;
          lut[5338] <= 16'd18732;
          lut[5339] <= 16'd18800;
          lut[5340] <= 16'd18867;
          lut[5341] <= 16'd18933;
          lut[5342] <= 16'd18997;
          lut[5343] <= 16'd19061;
          lut[5344] <= 16'd19123;
          lut[5345] <= 16'd19184;
          lut[5346] <= 16'd19244;
          lut[5347] <= 16'd19303;
          lut[5348] <= 16'd19361;
          lut[5349] <= 16'd19418;
          lut[5350] <= 16'd19474;
          lut[5351] <= 16'd19529;
          lut[5352] <= 16'd19583;
          lut[5353] <= 16'd19637;
          lut[5354] <= 16'd19689;
          lut[5355] <= 16'd19741;
          lut[5356] <= 16'd19791;
          lut[5357] <= 16'd19841;
          lut[5358] <= 16'd19890;
          lut[5359] <= 16'd19939;
          lut[5360] <= 16'd19986;
          lut[5361] <= 16'd20033;
          lut[5362] <= 16'd20079;
          lut[5363] <= 16'd20125;
          lut[5364] <= 16'd20170;
          lut[5365] <= 16'd20214;
          lut[5366] <= 16'd20257;
          lut[5367] <= 16'd20300;
          lut[5368] <= 16'd20342;
          lut[5369] <= 16'd20383;
          lut[5370] <= 16'd20424;
          lut[5371] <= 16'd20464;
          lut[5372] <= 16'd20504;
          lut[5373] <= 16'd20543;
          lut[5374] <= 16'd20582;
          lut[5375] <= 16'd20620;
          lut[5376] <= 0;
          lut[5377] <= 16'd390;
          lut[5378] <= 16'd780;
          lut[5379] <= 16'd1168;
          lut[5380] <= 16'd1556;
          lut[5381] <= 16'd1941;
          lut[5382] <= 16'd2325;
          lut[5383] <= 16'd2706;
          lut[5384] <= 16'd3084;
          lut[5385] <= 16'd3459;
          lut[5386] <= 16'd3830;
          lut[5387] <= 16'd4197;
          lut[5388] <= 16'd4560;
          lut[5389] <= 16'd4918;
          lut[5390] <= 16'd5272;
          lut[5391] <= 16'd5620;
          lut[5392] <= 16'd5963;
          lut[5393] <= 16'd6301;
          lut[5394] <= 16'd6634;
          lut[5395] <= 16'd6960;
          lut[5396] <= 16'd7281;
          lut[5397] <= 16'd7596;
          lut[5398] <= 16'd7905;
          lut[5399] <= 16'd8209;
          lut[5400] <= 16'd8506;
          lut[5401] <= 16'd8797;
          lut[5402] <= 16'd9082;
          lut[5403] <= 16'd9361;
          lut[5404] <= 16'd9634;
          lut[5405] <= 16'd9901;
          lut[5406] <= 16'd10162;
          lut[5407] <= 16'd10418;
          lut[5408] <= 16'd10667;
          lut[5409] <= 16'd10911;
          lut[5410] <= 16'd11150;
          lut[5411] <= 16'd11383;
          lut[5412] <= 16'd11610;
          lut[5413] <= 16'd11832;
          lut[5414] <= 16'd12049;
          lut[5415] <= 16'd12261;
          lut[5416] <= 16'd12468;
          lut[5417] <= 16'd12671;
          lut[5418] <= 16'd12868;
          lut[5419] <= 16'd13061;
          lut[5420] <= 16'd13249;
          lut[5421] <= 16'd13433;
          lut[5422] <= 16'd13612;
          lut[5423] <= 16'd13787;
          lut[5424] <= 16'd13959;
          lut[5425] <= 16'd14126;
          lut[5426] <= 16'd14289;
          lut[5427] <= 16'd14449;
          lut[5428] <= 16'd14604;
          lut[5429] <= 16'd14757;
          lut[5430] <= 16'd14905;
          lut[5431] <= 16'd15051;
          lut[5432] <= 16'd15193;
          lut[5433] <= 16'd15332;
          lut[5434] <= 16'd15467;
          lut[5435] <= 16'd15600;
          lut[5436] <= 16'd15730;
          lut[5437] <= 16'd15857;
          lut[5438] <= 16'd15981;
          lut[5439] <= 16'd16102;
          lut[5440] <= 16'd16221;
          lut[5441] <= 16'd16337;
          lut[5442] <= 16'd16451;
          lut[5443] <= 16'd16562;
          lut[5444] <= 16'd16671;
          lut[5445] <= 16'd16777;
          lut[5446] <= 16'd16882;
          lut[5447] <= 16'd16984;
          lut[5448] <= 16'd17084;
          lut[5449] <= 16'd17182;
          lut[5450] <= 16'd17278;
          lut[5451] <= 16'd17372;
          lut[5452] <= 16'd17464;
          lut[5453] <= 16'd17555;
          lut[5454] <= 16'd17643;
          lut[5455] <= 16'd17730;
          lut[5456] <= 16'd17815;
          lut[5457] <= 16'd17899;
          lut[5458] <= 16'd17980;
          lut[5459] <= 16'd18061;
          lut[5460] <= 16'd18140;
          lut[5461] <= 16'd18217;
          lut[5462] <= 16'd18293;
          lut[5463] <= 16'd18367;
          lut[5464] <= 16'd18440;
          lut[5465] <= 16'd18512;
          lut[5466] <= 16'd18582;
          lut[5467] <= 16'd18651;
          lut[5468] <= 16'd18719;
          lut[5469] <= 16'd18786;
          lut[5470] <= 16'd18851;
          lut[5471] <= 16'd18916;
          lut[5472] <= 16'd18979;
          lut[5473] <= 16'd19041;
          lut[5474] <= 16'd19102;
          lut[5475] <= 16'd19162;
          lut[5476] <= 16'd19221;
          lut[5477] <= 16'd19279;
          lut[5478] <= 16'd19336;
          lut[5479] <= 16'd19392;
          lut[5480] <= 16'd19447;
          lut[5481] <= 16'd19502;
          lut[5482] <= 16'd19555;
          lut[5483] <= 16'd19608;
          lut[5484] <= 16'd19659;
          lut[5485] <= 16'd19710;
          lut[5486] <= 16'd19760;
          lut[5487] <= 16'd19809;
          lut[5488] <= 16'd19858;
          lut[5489] <= 16'd19906;
          lut[5490] <= 16'd19953;
          lut[5491] <= 16'd19999;
          lut[5492] <= 16'd20044;
          lut[5493] <= 16'd20089;
          lut[5494] <= 16'd20133;
          lut[5495] <= 16'd20177;
          lut[5496] <= 16'd20220;
          lut[5497] <= 16'd20262;
          lut[5498] <= 16'd20304;
          lut[5499] <= 16'd20345;
          lut[5500] <= 16'd20385;
          lut[5501] <= 16'd20425;
          lut[5502] <= 16'd20464;
          lut[5503] <= 16'd20503;
          lut[5504] <= 0;
          lut[5505] <= 16'd381;
          lut[5506] <= 16'd761;
          lut[5507] <= 16'd1141;
          lut[5508] <= 16'd1520;
          lut[5509] <= 16'd1897;
          lut[5510] <= 16'd2271;
          lut[5511] <= 16'd2644;
          lut[5512] <= 16'd3014;
          lut[5513] <= 16'd3380;
          lut[5514] <= 16'd3744;
          lut[5515] <= 16'd4103;
          lut[5516] <= 16'd4459;
          lut[5517] <= 16'd4810;
          lut[5518] <= 16'd5157;
          lut[5519] <= 16'd5499;
          lut[5520] <= 16'd5836;
          lut[5521] <= 16'd6168;
          lut[5522] <= 16'd6495;
          lut[5523] <= 16'd6817;
          lut[5524] <= 16'd7133;
          lut[5525] <= 16'd7443;
          lut[5526] <= 16'd7748;
          lut[5527] <= 16'd8047;
          lut[5528] <= 16'd8341;
          lut[5529] <= 16'd8628;
          lut[5530] <= 16'd8910;
          lut[5531] <= 16'd9186;
          lut[5532] <= 16'd9457;
          lut[5533] <= 16'd9721;
          lut[5534] <= 16'd9981;
          lut[5535] <= 16'd10234;
          lut[5536] <= 16'd10482;
          lut[5537] <= 16'd10724;
          lut[5538] <= 16'd10962;
          lut[5539] <= 16'd11193;
          lut[5540] <= 16'd11420;
          lut[5541] <= 16'd11641;
          lut[5542] <= 16'd11858;
          lut[5543] <= 16'd12069;
          lut[5544] <= 16'd12276;
          lut[5545] <= 16'd12478;
          lut[5546] <= 16'd12675;
          lut[5547] <= 16'd12868;
          lut[5548] <= 16'd13056;
          lut[5549] <= 16'd13240;
          lut[5550] <= 16'd13420;
          lut[5551] <= 16'd13596;
          lut[5552] <= 16'd13767;
          lut[5553] <= 16'd13935;
          lut[5554] <= 16'd14099;
          lut[5555] <= 16'd14259;
          lut[5556] <= 16'd14416;
          lut[5557] <= 16'd14568;
          lut[5558] <= 16'd14718;
          lut[5559] <= 16'd14864;
          lut[5560] <= 16'd15007;
          lut[5561] <= 16'd15147;
          lut[5562] <= 16'd15284;
          lut[5563] <= 16'd15417;
          lut[5564] <= 16'd15548;
          lut[5565] <= 16'd15676;
          lut[5566] <= 16'd15801;
          lut[5567] <= 16'd15923;
          lut[5568] <= 16'd16043;
          lut[5569] <= 16'd16160;
          lut[5570] <= 16'd16275;
          lut[5571] <= 16'd16387;
          lut[5572] <= 16'd16497;
          lut[5573] <= 16'd16605;
          lut[5574] <= 16'd16711;
          lut[5575] <= 16'd16814;
          lut[5576] <= 16'd16915;
          lut[5577] <= 16'd17014;
          lut[5578] <= 16'd17112;
          lut[5579] <= 16'd17207;
          lut[5580] <= 16'd17300;
          lut[5581] <= 16'd17392;
          lut[5582] <= 16'd17481;
          lut[5583] <= 16'd17569;
          lut[5584] <= 16'd17655;
          lut[5585] <= 16'd17740;
          lut[5586] <= 16'd17823;
          lut[5587] <= 16'd17904;
          lut[5588] <= 16'd17984;
          lut[5589] <= 16'd18063;
          lut[5590] <= 16'd18140;
          lut[5591] <= 16'd18215;
          lut[5592] <= 16'd18289;
          lut[5593] <= 16'd18362;
          lut[5594] <= 16'd18433;
          lut[5595] <= 16'd18504;
          lut[5596] <= 16'd18572;
          lut[5597] <= 16'd18640;
          lut[5598] <= 16'd18707;
          lut[5599] <= 16'd18772;
          lut[5600] <= 16'd18836;
          lut[5601] <= 16'd18899;
          lut[5602] <= 16'd18961;
          lut[5603] <= 16'd19022;
          lut[5604] <= 16'd19082;
          lut[5605] <= 16'd19141;
          lut[5606] <= 16'd19199;
          lut[5607] <= 16'd19256;
          lut[5608] <= 16'd19312;
          lut[5609] <= 16'd19368;
          lut[5610] <= 16'd19422;
          lut[5611] <= 16'd19475;
          lut[5612] <= 16'd19528;
          lut[5613] <= 16'd19580;
          lut[5614] <= 16'd19631;
          lut[5615] <= 16'd19681;
          lut[5616] <= 16'd19730;
          lut[5617] <= 16'd19779;
          lut[5618] <= 16'd19826;
          lut[5619] <= 16'd19873;
          lut[5620] <= 16'd19920;
          lut[5621] <= 16'd19966;
          lut[5622] <= 16'd20011;
          lut[5623] <= 16'd20055;
          lut[5624] <= 16'd20099;
          lut[5625] <= 16'd20142;
          lut[5626] <= 16'd20184;
          lut[5627] <= 16'd20226;
          lut[5628] <= 16'd20267;
          lut[5629] <= 16'd20308;
          lut[5630] <= 16'd20348;
          lut[5631] <= 16'd20387;
          lut[5632] <= 0;
          lut[5633] <= 16'd372;
          lut[5634] <= 16'd744;
          lut[5635] <= 16'd1115;
          lut[5636] <= 16'd1485;
          lut[5637] <= 16'd1854;
          lut[5638] <= 16'd2220;
          lut[5639] <= 16'd2585;
          lut[5640] <= 16'd2947;
          lut[5641] <= 16'd3306;
          lut[5642] <= 16'd3661;
          lut[5643] <= 16'd4014;
          lut[5644] <= 16'd4362;
          lut[5645] <= 16'd4707;
          lut[5646] <= 16'd5047;
          lut[5647] <= 16'd5383;
          lut[5648] <= 16'd5714;
          lut[5649] <= 16'd6041;
          lut[5650] <= 16'd6362;
          lut[5651] <= 16'd6679;
          lut[5652] <= 16'd6990;
          lut[5653] <= 16'd7296;
          lut[5654] <= 16'd7596;
          lut[5655] <= 16'd7892;
          lut[5656] <= 16'd8181;
          lut[5657] <= 16'd8466;
          lut[5658] <= 16'd8744;
          lut[5659] <= 16'd9018;
          lut[5660] <= 16'd9285;
          lut[5661] <= 16'd9548;
          lut[5662] <= 16'd9804;
          lut[5663] <= 16'd10056;
          lut[5664] <= 16'd10302;
          lut[5665] <= 16'd10543;
          lut[5666] <= 16'd10779;
          lut[5667] <= 16'd11009;
          lut[5668] <= 16'd11235;
          lut[5669] <= 16'd11456;
          lut[5670] <= 16'd11671;
          lut[5671] <= 16'd11882;
          lut[5672] <= 16'd12088;
          lut[5673] <= 16'd12290;
          lut[5674] <= 16'd12487;
          lut[5675] <= 16'd12680;
          lut[5676] <= 16'd12868;
          lut[5677] <= 16'd13052;
          lut[5678] <= 16'd13232;
          lut[5679] <= 16'd13408;
          lut[5680] <= 16'd13580;
          lut[5681] <= 16'd13748;
          lut[5682] <= 16'd13912;
          lut[5683] <= 16'd14073;
          lut[5684] <= 16'd14230;
          lut[5685] <= 16'd14384;
          lut[5686] <= 16'd14534;
          lut[5687] <= 16'd14681;
          lut[5688] <= 16'd14825;
          lut[5689] <= 16'd14965;
          lut[5690] <= 16'd15103;
          lut[5691] <= 16'd15237;
          lut[5692] <= 16'd15369;
          lut[5693] <= 16'd15498;
          lut[5694] <= 16'd15624;
          lut[5695] <= 16'd15747;
          lut[5696] <= 16'd15868;
          lut[5697] <= 16'd15986;
          lut[5698] <= 16'd16102;
          lut[5699] <= 16'd16215;
          lut[5700] <= 16'd16327;
          lut[5701] <= 16'd16435;
          lut[5702] <= 16'd16542;
          lut[5703] <= 16'd16646;
          lut[5704] <= 16'd16748;
          lut[5705] <= 16'd16849;
          lut[5706] <= 16'd16947;
          lut[5707] <= 16'd17043;
          lut[5708] <= 16'd17138;
          lut[5709] <= 16'd17230;
          lut[5710] <= 16'd17321;
          lut[5711] <= 16'd17410;
          lut[5712] <= 16'd17497;
          lut[5713] <= 16'd17583;
          lut[5714] <= 16'd17667;
          lut[5715] <= 16'd17750;
          lut[5716] <= 16'd17830;
          lut[5717] <= 16'd17910;
          lut[5718] <= 16'd17988;
          lut[5719] <= 16'd18064;
          lut[5720] <= 16'd18140;
          lut[5721] <= 16'd18213;
          lut[5722] <= 16'd18286;
          lut[5723] <= 16'd18357;
          lut[5724] <= 16'd18427;
          lut[5725] <= 16'd18496;
          lut[5726] <= 16'd18563;
          lut[5727] <= 16'd18629;
          lut[5728] <= 16'd18695;
          lut[5729] <= 16'd18759;
          lut[5730] <= 16'd18822;
          lut[5731] <= 16'd18884;
          lut[5732] <= 16'd18945;
          lut[5733] <= 16'd19005;
          lut[5734] <= 16'd19063;
          lut[5735] <= 16'd19121;
          lut[5736] <= 16'd19178;
          lut[5737] <= 16'd19234;
          lut[5738] <= 16'd19290;
          lut[5739] <= 16'd19344;
          lut[5740] <= 16'd19397;
          lut[5741] <= 16'd19450;
          lut[5742] <= 16'd19502;
          lut[5743] <= 16'd19553;
          lut[5744] <= 16'd19603;
          lut[5745] <= 16'd19652;
          lut[5746] <= 16'd19701;
          lut[5747] <= 16'd19749;
          lut[5748] <= 16'd19796;
          lut[5749] <= 16'd19842;
          lut[5750] <= 16'd19888;
          lut[5751] <= 16'd19933;
          lut[5752] <= 16'd19978;
          lut[5753] <= 16'd20022;
          lut[5754] <= 16'd20065;
          lut[5755] <= 16'd20107;
          lut[5756] <= 16'd20149;
          lut[5757] <= 16'd20191;
          lut[5758] <= 16'd20231;
          lut[5759] <= 16'd20272;
          lut[5760] <= 0;
          lut[5761] <= 16'd364;
          lut[5762] <= 16'd728;
          lut[5763] <= 16'd1091;
          lut[5764] <= 16'd1453;
          lut[5765] <= 16'd1813;
          lut[5766] <= 16'd2172;
          lut[5767] <= 16'd2528;
          lut[5768] <= 16'd2883;
          lut[5769] <= 16'd3234;
          lut[5770] <= 16'd3583;
          lut[5771] <= 16'd3928;
          lut[5772] <= 16'd4270;
          lut[5773] <= 16'd4608;
          lut[5774] <= 16'd4942;
          lut[5775] <= 16'd5272;
          lut[5776] <= 16'd5597;
          lut[5777] <= 16'd5918;
          lut[5778] <= 16'd6234;
          lut[5779] <= 16'd6546;
          lut[5780] <= 16'd6852;
          lut[5781] <= 16'd7154;
          lut[5782] <= 16'd7450;
          lut[5783] <= 16'd7741;
          lut[5784] <= 16'd8027;
          lut[5785] <= 16'd8308;
          lut[5786] <= 16'd8584;
          lut[5787] <= 16'd8854;
          lut[5788] <= 16'd9119;
          lut[5789] <= 16'd9379;
          lut[5790] <= 16'd9634;
          lut[5791] <= 16'd9883;
          lut[5792] <= 16'd10128;
          lut[5793] <= 16'd10367;
          lut[5794] <= 16'd10601;
          lut[5795] <= 16'd10831;
          lut[5796] <= 16'd11055;
          lut[5797] <= 16'd11275;
          lut[5798] <= 16'd11489;
          lut[5799] <= 16'd11700;
          lut[5800] <= 16'd11905;
          lut[5801] <= 16'd12106;
          lut[5802] <= 16'd12303;
          lut[5803] <= 16'd12496;
          lut[5804] <= 16'd12684;
          lut[5805] <= 16'd12868;
          lut[5806] <= 16'd13048;
          lut[5807] <= 16'd13224;
          lut[5808] <= 16'd13396;
          lut[5809] <= 16'd13565;
          lut[5810] <= 16'd13729;
          lut[5811] <= 16'd13891;
          lut[5812] <= 16'd14048;
          lut[5813] <= 16'd14202;
          lut[5814] <= 16'd14353;
          lut[5815] <= 16'd14501;
          lut[5816] <= 16'd14645;
          lut[5817] <= 16'd14787;
          lut[5818] <= 16'd14925;
          lut[5819] <= 16'd15060;
          lut[5820] <= 16'd15193;
          lut[5821] <= 16'd15322;
          lut[5822] <= 16'd15449;
          lut[5823] <= 16'd15574;
          lut[5824] <= 16'd15695;
          lut[5825] <= 16'd15815;
          lut[5826] <= 16'd15931;
          lut[5827] <= 16'd16046;
          lut[5828] <= 16'd16158;
          lut[5829] <= 16'd16268;
          lut[5830] <= 16'd16375;
          lut[5831] <= 16'd16481;
          lut[5832] <= 16'd16584;
          lut[5833] <= 16'd16685;
          lut[5834] <= 16'd16784;
          lut[5835] <= 16'd16882;
          lut[5836] <= 16'd16977;
          lut[5837] <= 16'd17071;
          lut[5838] <= 16'd17163;
          lut[5839] <= 16'd17253;
          lut[5840] <= 16'd17341;
          lut[5841] <= 16'd17428;
          lut[5842] <= 16'd17513;
          lut[5843] <= 16'd17596;
          lut[5844] <= 16'd17678;
          lut[5845] <= 16'd17759;
          lut[5846] <= 16'd17838;
          lut[5847] <= 16'd17915;
          lut[5848] <= 16'd17991;
          lut[5849] <= 16'd18066;
          lut[5850] <= 16'd18140;
          lut[5851] <= 16'd18212;
          lut[5852] <= 16'd18283;
          lut[5853] <= 16'd18352;
          lut[5854] <= 16'd18421;
          lut[5855] <= 16'd18488;
          lut[5856] <= 16'd18554;
          lut[5857] <= 16'd18619;
          lut[5858] <= 16'd18683;
          lut[5859] <= 16'd18746;
          lut[5860] <= 16'd18808;
          lut[5861] <= 16'd18869;
          lut[5862] <= 16'd18929;
          lut[5863] <= 16'd18987;
          lut[5864] <= 16'd19045;
          lut[5865] <= 16'd19102;
          lut[5866] <= 16'd19158;
          lut[5867] <= 16'd19213;
          lut[5868] <= 16'd19268;
          lut[5869] <= 16'd19321;
          lut[5870] <= 16'd19374;
          lut[5871] <= 16'd19426;
          lut[5872] <= 16'd19477;
          lut[5873] <= 16'd19527;
          lut[5874] <= 16'd19576;
          lut[5875] <= 16'd19625;
          lut[5876] <= 16'd19673;
          lut[5877] <= 16'd19720;
          lut[5878] <= 16'd19767;
          lut[5879] <= 16'd19813;
          lut[5880] <= 16'd19858;
          lut[5881] <= 16'd19902;
          lut[5882] <= 16'd19946;
          lut[5883] <= 16'd19990;
          lut[5884] <= 16'd20032;
          lut[5885] <= 16'd20074;
          lut[5886] <= 16'd20116;
          lut[5887] <= 16'd20157;
          lut[5888] <= 0;
          lut[5889] <= 16'd356;
          lut[5890] <= 16'd712;
          lut[5891] <= 16'd1067;
          lut[5892] <= 16'd1421;
          lut[5893] <= 16'd1774;
          lut[5894] <= 16'd2125;
          lut[5895] <= 16'd2474;
          lut[5896] <= 16'd2821;
          lut[5897] <= 16'd3166;
          lut[5898] <= 16'd3507;
          lut[5899] <= 16'd3846;
          lut[5900] <= 16'd4181;
          lut[5901] <= 16'd4513;
          lut[5902] <= 16'd4841;
          lut[5903] <= 16'd5164;
          lut[5904] <= 16'd5484;
          lut[5905] <= 16'd5800;
          lut[5906] <= 16'd6111;
          lut[5907] <= 16'd6418;
          lut[5908] <= 16'd6720;
          lut[5909] <= 16'd7017;
          lut[5910] <= 16'd7309;
          lut[5911] <= 16'd7596;
          lut[5912] <= 16'd7879;
          lut[5913] <= 16'd8156;
          lut[5914] <= 16'd8429;
          lut[5915] <= 16'd8696;
          lut[5916] <= 16'd8959;
          lut[5917] <= 16'd9216;
          lut[5918] <= 16'd9468;
          lut[5919] <= 16'd9716;
          lut[5920] <= 16'd9958;
          lut[5921] <= 16'd10196;
          lut[5922] <= 16'd10429;
          lut[5923] <= 16'd10657;
          lut[5924] <= 16'd10880;
          lut[5925] <= 16'd11098;
          lut[5926] <= 16'd11312;
          lut[5927] <= 16'd11522;
          lut[5928] <= 16'd11727;
          lut[5929] <= 16'd11927;
          lut[5930] <= 16'd12124;
          lut[5931] <= 16'd12316;
          lut[5932] <= 16'd12504;
          lut[5933] <= 16'd12688;
          lut[5934] <= 16'd12868;
          lut[5935] <= 16'd13044;
          lut[5936] <= 16'd13217;
          lut[5937] <= 16'd13385;
          lut[5938] <= 16'd13550;
          lut[5939] <= 16'd13712;
          lut[5940] <= 16'd13870;
          lut[5941] <= 16'd14025;
          lut[5942] <= 16'd14176;
          lut[5943] <= 16'd14324;
          lut[5944] <= 16'd14469;
          lut[5945] <= 16'd14611;
          lut[5946] <= 16'd14750;
          lut[5947] <= 16'd14886;
          lut[5948] <= 16'd15019;
          lut[5949] <= 16'd15150;
          lut[5950] <= 16'd15278;
          lut[5951] <= 16'd15403;
          lut[5952] <= 16'd15525;
          lut[5953] <= 16'd15646;
          lut[5954] <= 16'd15763;
          lut[5955] <= 16'd15878;
          lut[5956] <= 16'd15991;
          lut[5957] <= 16'd16102;
          lut[5958] <= 16'd16211;
          lut[5959] <= 16'd16317;
          lut[5960] <= 16'd16421;
          lut[5961] <= 16'd16523;
          lut[5962] <= 16'd16624;
          lut[5963] <= 16'd16722;
          lut[5964] <= 16'd16818;
          lut[5965] <= 16'd16913;
          lut[5966] <= 16'd17006;
          lut[5967] <= 16'd17097;
          lut[5968] <= 16'd17186;
          lut[5969] <= 16'd17274;
          lut[5970] <= 16'd17360;
          lut[5971] <= 16'd17444;
          lut[5972] <= 16'd17527;
          lut[5973] <= 16'd17609;
          lut[5974] <= 16'd17689;
          lut[5975] <= 16'd17767;
          lut[5976] <= 16'd17844;
          lut[5977] <= 16'd17920;
          lut[5978] <= 16'd17995;
          lut[5979] <= 16'd18068;
          lut[5980] <= 16'd18140;
          lut[5981] <= 16'd18210;
          lut[5982] <= 16'd18280;
          lut[5983] <= 16'd18348;
          lut[5984] <= 16'd18415;
          lut[5985] <= 16'd18481;
          lut[5986] <= 16'd18546;
          lut[5987] <= 16'd18609;
          lut[5988] <= 16'd18672;
          lut[5989] <= 16'd18734;
          lut[5990] <= 16'd18795;
          lut[5991] <= 16'd18854;
          lut[5992] <= 16'd18913;
          lut[5993] <= 16'd18971;
          lut[5994] <= 16'd19028;
          lut[5995] <= 16'd19084;
          lut[5996] <= 16'd19139;
          lut[5997] <= 16'd19193;
          lut[5998] <= 16'd19247;
          lut[5999] <= 16'd19299;
          lut[6000] <= 16'd19351;
          lut[6001] <= 16'd19402;
          lut[6002] <= 16'd19452;
          lut[6003] <= 16'd19502;
          lut[6004] <= 16'd19550;
          lut[6005] <= 16'd19599;
          lut[6006] <= 16'd19646;
          lut[6007] <= 16'd19692;
          lut[6008] <= 16'd19738;
          lut[6009] <= 16'd19784;
          lut[6010] <= 16'd19828;
          lut[6011] <= 16'd19872;
          lut[6012] <= 16'd19916;
          lut[6013] <= 16'd19959;
          lut[6014] <= 16'd20001;
          lut[6015] <= 16'd20042;
          lut[6016] <= 0;
          lut[6017] <= 16'd349;
          lut[6018] <= 16'd697;
          lut[6019] <= 16'd1044;
          lut[6020] <= 16'd1391;
          lut[6021] <= 16'd1736;
          lut[6022] <= 16'd2080;
          lut[6023] <= 16'd2422;
          lut[6024] <= 16'd2762;
          lut[6025] <= 16'd3100;
          lut[6026] <= 16'd3435;
          lut[6027] <= 16'd3767;
          lut[6028] <= 16'd4096;
          lut[6029] <= 16'd4421;
          lut[6030] <= 16'd4743;
          lut[6031] <= 16'd5062;
          lut[6032] <= 16'd5376;
          lut[6033] <= 16'd5686;
          lut[6034] <= 16'd5992;
          lut[6035] <= 16'd6294;
          lut[6036] <= 16'd6592;
          lut[6037] <= 16'd6885;
          lut[6038] <= 16'd7173;
          lut[6039] <= 16'd7456;
          lut[6040] <= 16'd7735;
          lut[6041] <= 16'd8009;
          lut[6042] <= 16'd8279;
          lut[6043] <= 16'd8543;
          lut[6044] <= 16'd8803;
          lut[6045] <= 16'd9058;
          lut[6046] <= 16'd9308;
          lut[6047] <= 16'd9553;
          lut[6048] <= 16'd9794;
          lut[6049] <= 16'd10030;
          lut[6050] <= 16'd10261;
          lut[6051] <= 16'd10487;
          lut[6052] <= 16'd10709;
          lut[6053] <= 16'd10927;
          lut[6054] <= 16'd11140;
          lut[6055] <= 16'd11348;
          lut[6056] <= 16'd11553;
          lut[6057] <= 16'd11753;
          lut[6058] <= 16'd11948;
          lut[6059] <= 16'd12140;
          lut[6060] <= 16'd12328;
          lut[6061] <= 16'd12512;
          lut[6062] <= 16'd12692;
          lut[6063] <= 16'd12868;
          lut[6064] <= 16'd13040;
          lut[6065] <= 16'd13209;
          lut[6066] <= 16'd13375;
          lut[6067] <= 16'd13536;
          lut[6068] <= 16'd13695;
          lut[6069] <= 16'd13850;
          lut[6070] <= 16'd14002;
          lut[6071] <= 16'd14150;
          lut[6072] <= 16'd14296;
          lut[6073] <= 16'd14439;
          lut[6074] <= 16'd14578;
          lut[6075] <= 16'd14715;
          lut[6076] <= 16'd14849;
          lut[6077] <= 16'd14980;
          lut[6078] <= 16'd15109;
          lut[6079] <= 16'd15234;
          lut[6080] <= 16'd15358;
          lut[6081] <= 16'd15479;
          lut[6082] <= 16'd15597;
          lut[6083] <= 16'd15713;
          lut[6084] <= 16'd15827;
          lut[6085] <= 16'd15939;
          lut[6086] <= 16'd16048;
          lut[6087] <= 16'd16155;
          lut[6088] <= 16'd16261;
          lut[6089] <= 16'd16364;
          lut[6090] <= 16'd16465;
          lut[6091] <= 16'd16564;
          lut[6092] <= 16'd16662;
          lut[6093] <= 16'd16757;
          lut[6094] <= 16'd16851;
          lut[6095] <= 16'd16943;
          lut[6096] <= 16'd17033;
          lut[6097] <= 16'd17122;
          lut[6098] <= 16'd17209;
          lut[6099] <= 16'd17294;
          lut[6100] <= 16'd17378;
          lut[6101] <= 16'd17460;
          lut[6102] <= 16'd17541;
          lut[6103] <= 16'd17621;
          lut[6104] <= 16'd17699;
          lut[6105] <= 16'd17775;
          lut[6106] <= 16'd17851;
          lut[6107] <= 16'd17925;
          lut[6108] <= 16'd17998;
          lut[6109] <= 16'd18069;
          lut[6110] <= 16'd18140;
          lut[6111] <= 16'd18209;
          lut[6112] <= 16'd18277;
          lut[6113] <= 16'd18343;
          lut[6114] <= 16'd18409;
          lut[6115] <= 16'd18474;
          lut[6116] <= 16'd18537;
          lut[6117] <= 16'd18600;
          lut[6118] <= 16'd18662;
          lut[6119] <= 16'd18722;
          lut[6120] <= 16'd18782;
          lut[6121] <= 16'd18840;
          lut[6122] <= 16'd18898;
          lut[6123] <= 16'd18955;
          lut[6124] <= 16'd19011;
          lut[6125] <= 16'd19066;
          lut[6126] <= 16'd19120;
          lut[6127] <= 16'd19174;
          lut[6128] <= 16'd19226;
          lut[6129] <= 16'd19278;
          lut[6130] <= 16'd19329;
          lut[6131] <= 16'd19379;
          lut[6132] <= 16'd19429;
          lut[6133] <= 16'd19478;
          lut[6134] <= 16'd19526;
          lut[6135] <= 16'd19573;
          lut[6136] <= 16'd19620;
          lut[6137] <= 16'd19666;
          lut[6138] <= 16'd19711;
          lut[6139] <= 16'd19756;
          lut[6140] <= 16'd19800;
          lut[6141] <= 16'd19843;
          lut[6142] <= 16'd19886;
          lut[6143] <= 16'd19929;
          lut[6144] <= 0;
          lut[6145] <= 16'd341;
          lut[6146] <= 16'd682;
          lut[6147] <= 16'd1023;
          lut[6148] <= 16'd1362;
          lut[6149] <= 16'd1701;
          lut[6150] <= 16'd2037;
          lut[6151] <= 16'd2373;
          lut[6152] <= 16'd2706;
          lut[6153] <= 16'd3037;
          lut[6154] <= 16'd3365;
          lut[6155] <= 16'd3691;
          lut[6156] <= 16'd4014;
          lut[6157] <= 16'd4333;
          lut[6158] <= 16'd4650;
          lut[6159] <= 16'd4962;
          lut[6160] <= 16'd5272;
          lut[6161] <= 16'd5577;
          lut[6162] <= 16'd5878;
          lut[6163] <= 16'd6175;
          lut[6164] <= 16'd6468;
          lut[6165] <= 16'd6757;
          lut[6166] <= 16'd7041;
          lut[6167] <= 16'd7321;
          lut[6168] <= 16'd7596;
          lut[6169] <= 16'd7867;
          lut[6170] <= 16'd8133;
          lut[6171] <= 16'd8395;
          lut[6172] <= 16'd8652;
          lut[6173] <= 16'd8904;
          lut[6174] <= 16'd9152;
          lut[6175] <= 16'd9395;
          lut[6176] <= 16'd9634;
          lut[6177] <= 16'd9868;
          lut[6178] <= 16'd10097;
          lut[6179] <= 16'd10322;
          lut[6180] <= 16'd10543;
          lut[6181] <= 16'd10759;
          lut[6182] <= 16'd10971;
          lut[6183] <= 16'd11179;
          lut[6184] <= 16'd11383;
          lut[6185] <= 16'd11582;
          lut[6186] <= 16'd11777;
          lut[6187] <= 16'd11969;
          lut[6188] <= 16'd12156;
          lut[6189] <= 16'd12340;
          lut[6190] <= 16'd12519;
          lut[6191] <= 16'd12696;
          lut[6192] <= 16'd12868;
          lut[6193] <= 16'd13037;
          lut[6194] <= 16'd13202;
          lut[6195] <= 16'd13364;
          lut[6196] <= 16'd13523;
          lut[6197] <= 16'd13678;
          lut[6198] <= 16'd13831;
          lut[6199] <= 16'd13980;
          lut[6200] <= 16'd14126;
          lut[6201] <= 16'd14269;
          lut[6202] <= 16'd14409;
          lut[6203] <= 16'd14546;
          lut[6204] <= 16'd14681;
          lut[6205] <= 16'd14813;
          lut[6206] <= 16'd14942;
          lut[6207] <= 16'd15069;
          lut[6208] <= 16'd15193;
          lut[6209] <= 16'd15314;
          lut[6210] <= 16'd15434;
          lut[6211] <= 16'd15551;
          lut[6212] <= 16'd15665;
          lut[6213] <= 16'd15778;
          lut[6214] <= 16'd15888;
          lut[6215] <= 16'd15996;
          lut[6216] <= 16'd16102;
          lut[6217] <= 16'd16206;
          lut[6218] <= 16'd16308;
          lut[6219] <= 16'd16408;
          lut[6220] <= 16'd16507;
          lut[6221] <= 16'd16603;
          lut[6222] <= 16'd16698;
          lut[6223] <= 16'd16791;
          lut[6224] <= 16'd16882;
          lut[6225] <= 16'd16971;
          lut[6226] <= 16'd17059;
          lut[6227] <= 16'd17145;
          lut[6228] <= 16'd17230;
          lut[6229] <= 16'd17314;
          lut[6230] <= 16'd17395;
          lut[6231] <= 16'd17476;
          lut[6232] <= 16'd17555;
          lut[6233] <= 16'd17632;
          lut[6234] <= 16'd17708;
          lut[6235] <= 16'd17783;
          lut[6236] <= 16'd17857;
          lut[6237] <= 16'd17929;
          lut[6238] <= 16'd18001;
          lut[6239] <= 16'd18071;
          lut[6240] <= 16'd18140;
          lut[6241] <= 16'd18207;
          lut[6242] <= 16'd18274;
          lut[6243] <= 16'd18339;
          lut[6244] <= 16'd18404;
          lut[6245] <= 16'd18467;
          lut[6246] <= 16'd18530;
          lut[6247] <= 16'd18591;
          lut[6248] <= 16'd18651;
          lut[6249] <= 16'd18711;
          lut[6250] <= 16'd18769;
          lut[6251] <= 16'd18827;
          lut[6252] <= 16'd18884;
          lut[6253] <= 16'd18940;
          lut[6254] <= 16'd18995;
          lut[6255] <= 16'd19049;
          lut[6256] <= 16'd19102;
          lut[6257] <= 16'd19155;
          lut[6258] <= 16'd19207;
          lut[6259] <= 16'd19258;
          lut[6260] <= 16'd19308;
          lut[6261] <= 16'd19357;
          lut[6262] <= 16'd19406;
          lut[6263] <= 16'd19454;
          lut[6264] <= 16'd19502;
          lut[6265] <= 16'd19548;
          lut[6266] <= 16'd19595;
          lut[6267] <= 16'd19640;
          lut[6268] <= 16'd19685;
          lut[6269] <= 16'd19729;
          lut[6270] <= 16'd19772;
          lut[6271] <= 16'd19815;
          lut[6272] <= 0;
          lut[6273] <= 16'd334;
          lut[6274] <= 16'd668;
          lut[6275] <= 16'd1002;
          lut[6276] <= 16'd1335;
          lut[6277] <= 16'd1666;
          lut[6278] <= 16'd1996;
          lut[6279] <= 16'd2325;
          lut[6280] <= 16'd2652;
          lut[6281] <= 16'd2976;
          lut[6282] <= 16'd3298;
          lut[6283] <= 16'd3618;
          lut[6284] <= 16'd3935;
          lut[6285] <= 16'd4249;
          lut[6286] <= 16'd4560;
          lut[6287] <= 16'd4867;
          lut[6288] <= 16'd5171;
          lut[6289] <= 16'd5471;
          lut[6290] <= 16'd5768;
          lut[6291] <= 16'd6061;
          lut[6292] <= 16'd6349;
          lut[6293] <= 16'd6634;
          lut[6294] <= 16'd6914;
          lut[6295] <= 16'd7190;
          lut[6296] <= 16'd7462;
          lut[6297] <= 16'd7730;
          lut[6298] <= 16'd7993;
          lut[6299] <= 16'd8251;
          lut[6300] <= 16'd8506;
          lut[6301] <= 16'd8756;
          lut[6302] <= 16'd9001;
          lut[6303] <= 16'd9242;
          lut[6304] <= 16'd9479;
          lut[6305] <= 16'd9711;
          lut[6306] <= 16'd9939;
          lut[6307] <= 16'd10162;
          lut[6308] <= 16'd10381;
          lut[6309] <= 16'd10596;
          lut[6310] <= 16'd10807;
          lut[6311] <= 16'd11014;
          lut[6312] <= 16'd11217;
          lut[6313] <= 16'd11415;
          lut[6314] <= 16'd11610;
          lut[6315] <= 16'd11801;
          lut[6316] <= 16'd11988;
          lut[6317] <= 16'd12171;
          lut[6318] <= 16'd12351;
          lut[6319] <= 16'd12527;
          lut[6320] <= 16'd12699;
          lut[6321] <= 16'd12868;
          lut[6322] <= 16'd13033;
          lut[6323] <= 16'd13196;
          lut[6324] <= 16'd13354;
          lut[6325] <= 16'd13510;
          lut[6326] <= 16'd13663;
          lut[6327] <= 16'd13812;
          lut[6328] <= 16'd13959;
          lut[6329] <= 16'd14102;
          lut[6330] <= 16'd14243;
          lut[6331] <= 16'd14381;
          lut[6332] <= 16'd14516;
          lut[6333] <= 16'd14648;
          lut[6334] <= 16'd14778;
          lut[6335] <= 16'd14905;
          lut[6336] <= 16'd15030;
          lut[6337] <= 16'd15153;
          lut[6338] <= 16'd15273;
          lut[6339] <= 16'd15390;
          lut[6340] <= 16'd15506;
          lut[6341] <= 16'd15619;
          lut[6342] <= 16'd15730;
          lut[6343] <= 16'd15839;
          lut[6344] <= 16'd15946;
          lut[6345] <= 16'd16050;
          lut[6346] <= 16'd16153;
          lut[6347] <= 16'd16254;
          lut[6348] <= 16'd16353;
          lut[6349] <= 16'd16451;
          lut[6350] <= 16'd16546;
          lut[6351] <= 16'd16640;
          lut[6352] <= 16'd16732;
          lut[6353] <= 16'd16822;
          lut[6354] <= 16'd16911;
          lut[6355] <= 16'd16998;
          lut[6356] <= 16'd17084;
          lut[6357] <= 16'd17168;
          lut[6358] <= 16'd17251;
          lut[6359] <= 16'd17332;
          lut[6360] <= 16'd17412;
          lut[6361] <= 16'd17490;
          lut[6362] <= 16'd17567;
          lut[6363] <= 16'd17643;
          lut[6364] <= 16'd17718;
          lut[6365] <= 16'd17791;
          lut[6366] <= 16'd17863;
          lut[6367] <= 16'd17934;
          lut[6368] <= 16'd18004;
          lut[6369] <= 16'd18072;
          lut[6370] <= 16'd18140;
          lut[6371] <= 16'd18206;
          lut[6372] <= 16'd18271;
          lut[6373] <= 16'd18335;
          lut[6374] <= 16'd18399;
          lut[6375] <= 16'd18461;
          lut[6376] <= 16'd18522;
          lut[6377] <= 16'd18582;
          lut[6378] <= 16'd18642;
          lut[6379] <= 16'd18700;
          lut[6380] <= 16'd18757;
          lut[6381] <= 16'd18814;
          lut[6382] <= 16'd18870;
          lut[6383] <= 16'd18925;
          lut[6384] <= 16'd18979;
          lut[6385] <= 16'd19032;
          lut[6386] <= 16'd19085;
          lut[6387] <= 16'd19137;
          lut[6388] <= 16'd19188;
          lut[6389] <= 16'd19238;
          lut[6390] <= 16'd19287;
          lut[6391] <= 16'd19336;
          lut[6392] <= 16'd19384;
          lut[6393] <= 16'd19432;
          lut[6394] <= 16'd19479;
          lut[6395] <= 16'd19525;
          lut[6396] <= 16'd19570;
          lut[6397] <= 16'd19615;
          lut[6398] <= 16'd19659;
          lut[6399] <= 16'd19703;
          lut[6400] <= 0;
          lut[6401] <= 16'd328;
          lut[6402] <= 16'd655;
          lut[6403] <= 16'd982;
          lut[6404] <= 16'd1308;
          lut[6405] <= 16'd1633;
          lut[6406] <= 16'd1957;
          lut[6407] <= 16'd2279;
          lut[6408] <= 16'd2599;
          lut[6409] <= 16'd2918;
          lut[6410] <= 16'd3234;
          lut[6411] <= 16'd3548;
          lut[6412] <= 16'd3859;
          lut[6413] <= 16'd4168;
          lut[6414] <= 16'd4473;
          lut[6415] <= 16'd4775;
          lut[6416] <= 16'd5074;
          lut[6417] <= 16'd5370;
          lut[6418] <= 16'd5662;
          lut[6419] <= 16'd5950;
          lut[6420] <= 16'd6234;
          lut[6421] <= 16'd6515;
          lut[6422] <= 16'd6791;
          lut[6423] <= 16'd7064;
          lut[6424] <= 16'd7332;
          lut[6425] <= 16'd7596;
          lut[6426] <= 16'd7856;
          lut[6427] <= 16'd8112;
          lut[6428] <= 16'd8364;
          lut[6429] <= 16'd8611;
          lut[6430] <= 16'd8854;
          lut[6431] <= 16'd9093;
          lut[6432] <= 16'd9328;
          lut[6433] <= 16'd9558;
          lut[6434] <= 16'd9784;
          lut[6435] <= 16'd10006;
          lut[6436] <= 16'd10224;
          lut[6437] <= 16'd10438;
          lut[6438] <= 16'd10647;
          lut[6439] <= 16'd10853;
          lut[6440] <= 16'd11055;
          lut[6441] <= 16'd11253;
          lut[6442] <= 16'd11447;
          lut[6443] <= 16'd11637;
          lut[6444] <= 16'd11824;
          lut[6445] <= 16'd12006;
          lut[6446] <= 16'd12186;
          lut[6447] <= 16'd12361;
          lut[6448] <= 16'd12534;
          lut[6449] <= 16'd12702;
          lut[6450] <= 16'd12868;
          lut[6451] <= 16'd13030;
          lut[6452] <= 16'd13189;
          lut[6453] <= 16'd13345;
          lut[6454] <= 16'd13498;
          lut[6455] <= 16'd13648;
          lut[6456] <= 16'd13794;
          lut[6457] <= 16'd13938;
          lut[6458] <= 16'd14079;
          lut[6459] <= 16'd14218;
          lut[6460] <= 16'd14353;
          lut[6461] <= 16'd14486;
          lut[6462] <= 16'd14617;
          lut[6463] <= 16'd14745;
          lut[6464] <= 16'd14870;
          lut[6465] <= 16'd14993;
          lut[6466] <= 16'd15114;
          lut[6467] <= 16'd15232;
          lut[6468] <= 16'd15348;
          lut[6469] <= 16'd15462;
          lut[6470] <= 16'd15574;
          lut[6471] <= 16'd15683;
          lut[6472] <= 16'd15791;
          lut[6473] <= 16'd15897;
          lut[6474] <= 16'd16000;
          lut[6475] <= 16'd16102;
          lut[6476] <= 16'd16202;
          lut[6477] <= 16'd16300;
          lut[6478] <= 16'd16396;
          lut[6479] <= 16'd16491;
          lut[6480] <= 16'd16584;
          lut[6481] <= 16'd16675;
          lut[6482] <= 16'd16765;
          lut[6483] <= 16'd16853;
          lut[6484] <= 16'd16939;
          lut[6485] <= 16'd17024;
          lut[6486] <= 16'd17108;
          lut[6487] <= 16'd17190;
          lut[6488] <= 16'd17270;
          lut[6489] <= 16'd17350;
          lut[6490] <= 16'd17428;
          lut[6491] <= 16'd17504;
          lut[6492] <= 16'd17580;
          lut[6493] <= 16'd17654;
          lut[6494] <= 16'd17727;
          lut[6495] <= 16'd17798;
          lut[6496] <= 16'd17869;
          lut[6497] <= 16'd17938;
          lut[6498] <= 16'd18006;
          lut[6499] <= 16'd18073;
          lut[6500] <= 16'd18140;
          lut[6501] <= 16'd18205;
          lut[6502] <= 16'd18269;
          lut[6503] <= 16'd18332;
          lut[6504] <= 16'd18394;
          lut[6505] <= 16'd18455;
          lut[6506] <= 16'd18515;
          lut[6507] <= 16'd18574;
          lut[6508] <= 16'd18632;
          lut[6509] <= 16'd18690;
          lut[6510] <= 16'd18746;
          lut[6511] <= 16'd18802;
          lut[6512] <= 16'd18857;
          lut[6513] <= 16'd18911;
          lut[6514] <= 16'd18964;
          lut[6515] <= 16'd19016;
          lut[6516] <= 16'd19068;
          lut[6517] <= 16'd19119;
          lut[6518] <= 16'd19169;
          lut[6519] <= 16'd19219;
          lut[6520] <= 16'd19268;
          lut[6521] <= 16'd19316;
          lut[6522] <= 16'd19363;
          lut[6523] <= 16'd19410;
          lut[6524] <= 16'd19456;
          lut[6525] <= 16'd19502;
          lut[6526] <= 16'd19547;
          lut[6527] <= 16'd19591;
          lut[6528] <= 0;
          lut[6529] <= 16'd321;
          lut[6530] <= 16'd642;
          lut[6531] <= 16'd963;
          lut[6532] <= 16'd1282;
          lut[6533] <= 16'd1601;
          lut[6534] <= 16'd1919;
          lut[6535] <= 16'd2235;
          lut[6536] <= 16'd2549;
          lut[6537] <= 16'd2862;
          lut[6538] <= 16'd3172;
          lut[6539] <= 16'd3480;
          lut[6540] <= 16'd3786;
          lut[6541] <= 16'd4089;
          lut[6542] <= 16'd4389;
          lut[6543] <= 16'd4687;
          lut[6544] <= 16'd4981;
          lut[6545] <= 16'd5272;
          lut[6546] <= 16'd5559;
          lut[6547] <= 16'd5843;
          lut[6548] <= 16'd6123;
          lut[6549] <= 16'd6400;
          lut[6550] <= 16'd6672;
          lut[6551] <= 16'd6941;
          lut[6552] <= 16'd7206;
          lut[6553] <= 16'd7467;
          lut[6554] <= 16'd7724;
          lut[6555] <= 16'd7977;
          lut[6556] <= 16'd8226;
          lut[6557] <= 16'd8471;
          lut[6558] <= 16'd8712;
          lut[6559] <= 16'd8948;
          lut[6560] <= 16'd9181;
          lut[6561] <= 16'd9409;
          lut[6562] <= 16'd9634;
          lut[6563] <= 16'd9854;
          lut[6564] <= 16'd10071;
          lut[6565] <= 16'd10283;
          lut[6566] <= 16'd10492;
          lut[6567] <= 16'd10696;
          lut[6568] <= 16'd10897;
          lut[6569] <= 16'd11094;
          lut[6570] <= 16'd11287;
          lut[6571] <= 16'd11477;
          lut[6572] <= 16'd11663;
          lut[6573] <= 16'd11845;
          lut[6574] <= 16'd12024;
          lut[6575] <= 16'd12200;
          lut[6576] <= 16'd12372;
          lut[6577] <= 16'd12540;
          lut[6578] <= 16'd12706;
          lut[6579] <= 16'd12868;
          lut[6580] <= 16'd13027;
          lut[6581] <= 16'd13183;
          lut[6582] <= 16'd13336;
          lut[6583] <= 16'd13486;
          lut[6584] <= 16'd13633;
          lut[6585] <= 16'd13777;
          lut[6586] <= 16'd13919;
          lut[6587] <= 16'd14057;
          lut[6588] <= 16'd14193;
          lut[6589] <= 16'd14327;
          lut[6590] <= 16'd14458;
          lut[6591] <= 16'd14586;
          lut[6592] <= 16'd14712;
          lut[6593] <= 16'd14836;
          lut[6594] <= 16'd14957;
          lut[6595] <= 16'd15076;
          lut[6596] <= 16'd15193;
          lut[6597] <= 16'd15307;
          lut[6598] <= 16'd15420;
          lut[6599] <= 16'd15530;
          lut[6600] <= 16'd15639;
          lut[6601] <= 16'd15745;
          lut[6602] <= 16'd15849;
          lut[6603] <= 16'd15952;
          lut[6604] <= 16'd16052;
          lut[6605] <= 16'd16151;
          lut[6606] <= 16'd16248;
          lut[6607] <= 16'd16344;
          lut[6608] <= 16'd16437;
          lut[6609] <= 16'd16529;
          lut[6610] <= 16'd16620;
          lut[6611] <= 16'd16709;
          lut[6612] <= 16'd16796;
          lut[6613] <= 16'd16882;
          lut[6614] <= 16'd16966;
          lut[6615] <= 16'd17049;
          lut[6616] <= 16'd17130;
          lut[6617] <= 16'd17210;
          lut[6618] <= 16'd17289;
          lut[6619] <= 16'd17367;
          lut[6620] <= 16'd17443;
          lut[6621] <= 16'd17518;
          lut[6622] <= 16'd17591;
          lut[6623] <= 16'd17664;
          lut[6624] <= 16'd17735;
          lut[6625] <= 16'd17805;
          lut[6626] <= 16'd17874;
          lut[6627] <= 16'd17942;
          lut[6628] <= 16'd18009;
          lut[6629] <= 16'd18075;
          lut[6630] <= 16'd18140;
          lut[6631] <= 16'd18203;
          lut[6632] <= 16'd18266;
          lut[6633] <= 16'd18328;
          lut[6634] <= 16'd18389;
          lut[6635] <= 16'd18449;
          lut[6636] <= 16'd18508;
          lut[6637] <= 16'd18566;
          lut[6638] <= 16'd18623;
          lut[6639] <= 16'd18679;
          lut[6640] <= 16'd18735;
          lut[6641] <= 16'd18790;
          lut[6642] <= 16'd18844;
          lut[6643] <= 16'd18897;
          lut[6644] <= 16'd18949;
          lut[6645] <= 16'd19001;
          lut[6646] <= 16'd19052;
          lut[6647] <= 16'd19102;
          lut[6648] <= 16'd19152;
          lut[6649] <= 16'd19200;
          lut[6650] <= 16'd19249;
          lut[6651] <= 16'd19296;
          lut[6652] <= 16'd19343;
          lut[6653] <= 16'd19389;
          lut[6654] <= 16'd19435;
          lut[6655] <= 16'd19479;
          lut[6656] <= 0;
          lut[6657] <= 16'd315;
          lut[6658] <= 16'd630;
          lut[6659] <= 16'd944;
          lut[6660] <= 16'd1258;
          lut[6661] <= 16'd1571;
          lut[6662] <= 16'd1882;
          lut[6663] <= 16'd2192;
          lut[6664] <= 16'd2501;
          lut[6665] <= 16'd2808;
          lut[6666] <= 16'd3113;
          lut[6667] <= 16'd3415;
          lut[6668] <= 16'd3716;
          lut[6669] <= 16'd4014;
          lut[6670] <= 16'd4309;
          lut[6671] <= 16'd4601;
          lut[6672] <= 16'd4891;
          lut[6673] <= 16'd5177;
          lut[6674] <= 16'd5460;
          lut[6675] <= 16'd5740;
          lut[6676] <= 16'd6016;
          lut[6677] <= 16'd6288;
          lut[6678] <= 16'd6558;
          lut[6679] <= 16'd6823;
          lut[6680] <= 16'd7085;
          lut[6681] <= 16'd7342;
          lut[6682] <= 16'd7596;
          lut[6683] <= 16'd7847;
          lut[6684] <= 16'd8093;
          lut[6685] <= 16'd8335;
          lut[6686] <= 16'd8573;
          lut[6687] <= 16'd8808;
          lut[6688] <= 16'd9038;
          lut[6689] <= 16'd9265;
          lut[6690] <= 16'd9488;
          lut[6691] <= 16'd9706;
          lut[6692] <= 16'd9921;
          lut[6693] <= 16'd10132;
          lut[6694] <= 16'd10340;
          lut[6695] <= 16'd10543;
          lut[6696] <= 16'd10743;
          lut[6697] <= 16'd10939;
          lut[6698] <= 16'd11132;
          lut[6699] <= 16'd11320;
          lut[6700] <= 16'd11506;
          lut[6701] <= 16'd11688;
          lut[6702] <= 16'd11866;
          lut[6703] <= 16'd12041;
          lut[6704] <= 16'd12213;
          lut[6705] <= 16'd12381;
          lut[6706] <= 16'd12547;
          lut[6707] <= 16'd12709;
          lut[6708] <= 16'd12868;
          lut[6709] <= 16'd13024;
          lut[6710] <= 16'd13177;
          lut[6711] <= 16'd13327;
          lut[6712] <= 16'd13475;
          lut[6713] <= 16'd13619;
          lut[6714] <= 16'd13761;
          lut[6715] <= 16'd13900;
          lut[6716] <= 16'd14036;
          lut[6717] <= 16'd14170;
          lut[6718] <= 16'd14301;
          lut[6719] <= 16'd14430;
          lut[6720] <= 16'd14557;
          lut[6721] <= 16'd14681;
          lut[6722] <= 16'd14803;
          lut[6723] <= 16'd14922;
          lut[6724] <= 16'd15040;
          lut[6725] <= 16'd15155;
          lut[6726] <= 16'd15268;
          lut[6727] <= 16'd15379;
          lut[6728] <= 16'd15488;
          lut[6729] <= 16'd15595;
          lut[6730] <= 16'd15700;
          lut[6731] <= 16'd15803;
          lut[6732] <= 16'd15905;
          lut[6733] <= 16'd16004;
          lut[6734] <= 16'd16102;
          lut[6735] <= 16'd16198;
          lut[6736] <= 16'd16293;
          lut[6737] <= 16'd16385;
          lut[6738] <= 16'd16477;
          lut[6739] <= 16'd16566;
          lut[6740] <= 16'd16654;
          lut[6741] <= 16'd16741;
          lut[6742] <= 16'd16826;
          lut[6743] <= 16'd16909;
          lut[6744] <= 16'd16992;
          lut[6745] <= 16'd17073;
          lut[6746] <= 16'd17152;
          lut[6747] <= 16'd17230;
          lut[6748] <= 16'd17307;
          lut[6749] <= 16'd17383;
          lut[6750] <= 16'd17457;
          lut[6751] <= 16'd17530;
          lut[6752] <= 16'd17603;
          lut[6753] <= 16'd17673;
          lut[6754] <= 16'd17743;
          lut[6755] <= 16'd17812;
          lut[6756] <= 16'd17879;
          lut[6757] <= 16'd17946;
          lut[6758] <= 16'd18012;
          lut[6759] <= 16'd18076;
          lut[6760] <= 16'd18140;
          lut[6761] <= 16'd18202;
          lut[6762] <= 16'd18264;
          lut[6763] <= 16'd18324;
          lut[6764] <= 16'd18384;
          lut[6765] <= 16'd18443;
          lut[6766] <= 16'd18501;
          lut[6767] <= 16'd18558;
          lut[6768] <= 16'd18614;
          lut[6769] <= 16'd18670;
          lut[6770] <= 16'd18724;
          lut[6771] <= 16'd18778;
          lut[6772] <= 16'd18831;
          lut[6773] <= 16'd18884;
          lut[6774] <= 16'd18935;
          lut[6775] <= 16'd18986;
          lut[6776] <= 16'd19036;
          lut[6777] <= 16'd19086;
          lut[6778] <= 16'd19135;
          lut[6779] <= 16'd19183;
          lut[6780] <= 16'd19230;
          lut[6781] <= 16'd19277;
          lut[6782] <= 16'd19323;
          lut[6783] <= 16'd19369;
          lut[6784] <= 0;
          lut[6785] <= 16'd309;
          lut[6786] <= 16'd618;
          lut[6787] <= 16'd926;
          lut[6788] <= 16'd1234;
          lut[6789] <= 16'd1541;
          lut[6790] <= 16'd1847;
          lut[6791] <= 16'd2151;
          lut[6792] <= 16'd2455;
          lut[6793] <= 16'd2756;
          lut[6794] <= 16'd3055;
          lut[6795] <= 16'd3353;
          lut[6796] <= 16'd3648;
          lut[6797] <= 16'd3941;
          lut[6798] <= 16'd4231;
          lut[6799] <= 16'd4519;
          lut[6800] <= 16'd4804;
          lut[6801] <= 16'd5085;
          lut[6802] <= 16'd5364;
          lut[6803] <= 16'd5640;
          lut[6804] <= 16'd5912;
          lut[6805] <= 16'd6181;
          lut[6806] <= 16'd6446;
          lut[6807] <= 16'd6708;
          lut[6808] <= 16'd6967;
          lut[6809] <= 16'd7221;
          lut[6810] <= 16'd7472;
          lut[6811] <= 16'd7720;
          lut[6812] <= 16'd7963;
          lut[6813] <= 16'd8203;
          lut[6814] <= 16'd8439;
          lut[6815] <= 16'd8671;
          lut[6816] <= 16'd8900;
          lut[6817] <= 16'd9124;
          lut[6818] <= 16'd9345;
          lut[6819] <= 16'd9562;
          lut[6820] <= 16'd9776;
          lut[6821] <= 16'd9985;
          lut[6822] <= 16'd10191;
          lut[6823] <= 16'd10394;
          lut[6824] <= 16'd10592;
          lut[6825] <= 16'd10788;
          lut[6826] <= 16'd10979;
          lut[6827] <= 16'd11167;
          lut[6828] <= 16'd11352;
          lut[6829] <= 16'd11533;
          lut[6830] <= 16'd11711;
          lut[6831] <= 16'd11886;
          lut[6832] <= 16'd12058;
          lut[6833] <= 16'd12226;
          lut[6834] <= 16'd12391;
          lut[6835] <= 16'd12553;
          lut[6836] <= 16'd12712;
          lut[6837] <= 16'd12868;
          lut[6838] <= 16'd13021;
          lut[6839] <= 16'd13171;
          lut[6840] <= 16'd13319;
          lut[6841] <= 16'd13463;
          lut[6842] <= 16'd13605;
          lut[6843] <= 16'd13745;
          lut[6844] <= 16'd13882;
          lut[6845] <= 16'd14016;
          lut[6846] <= 16'd14148;
          lut[6847] <= 16'd14277;
          lut[6848] <= 16'd14404;
          lut[6849] <= 16'd14528;
          lut[6850] <= 16'd14651;
          lut[6851] <= 16'd14771;
          lut[6852] <= 16'd14889;
          lut[6853] <= 16'd15004;
          lut[6854] <= 16'd15118;
          lut[6855] <= 16'd15230;
          lut[6856] <= 16'd15339;
          lut[6857] <= 16'd15447;
          lut[6858] <= 16'd15553;
          lut[6859] <= 16'd15657;
          lut[6860] <= 16'd15759;
          lut[6861] <= 16'd15859;
          lut[6862] <= 16'd15958;
          lut[6863] <= 16'd16054;
          lut[6864] <= 16'd16149;
          lut[6865] <= 16'd16243;
          lut[6866] <= 16'd16335;
          lut[6867] <= 16'd16425;
          lut[6868] <= 16'd16514;
          lut[6869] <= 16'd16601;
          lut[6870] <= 16'd16687;
          lut[6871] <= 16'd16771;
          lut[6872] <= 16'd16854;
          lut[6873] <= 16'd16936;
          lut[6874] <= 16'd17016;
          lut[6875] <= 16'd17095;
          lut[6876] <= 16'd17173;
          lut[6877] <= 16'd17249;
          lut[6878] <= 16'd17324;
          lut[6879] <= 16'd17398;
          lut[6880] <= 16'd17471;
          lut[6881] <= 16'd17543;
          lut[6882] <= 16'd17613;
          lut[6883] <= 16'd17683;
          lut[6884] <= 16'd17751;
          lut[6885] <= 16'd17818;
          lut[6886] <= 16'd17885;
          lut[6887] <= 16'd17950;
          lut[6888] <= 16'd18014;
          lut[6889] <= 16'd18077;
          lut[6890] <= 16'd18140;
          lut[6891] <= 16'd18201;
          lut[6892] <= 16'd18261;
          lut[6893] <= 16'd18321;
          lut[6894] <= 16'd18380;
          lut[6895] <= 16'd18437;
          lut[6896] <= 16'd18494;
          lut[6897] <= 16'd18551;
          lut[6898] <= 16'd18606;
          lut[6899] <= 16'd18660;
          lut[6900] <= 16'd18714;
          lut[6901] <= 16'd18767;
          lut[6902] <= 16'd18819;
          lut[6903] <= 16'd18871;
          lut[6904] <= 16'd18922;
          lut[6905] <= 16'd18972;
          lut[6906] <= 16'd19021;
          lut[6907] <= 16'd19070;
          lut[6908] <= 16'd19118;
          lut[6909] <= 16'd19166;
          lut[6910] <= 16'd19212;
          lut[6911] <= 16'd19259;
          lut[6912] <= 0;
          lut[6913] <= 16'd303;
          lut[6914] <= 16'd607;
          lut[6915] <= 16'd909;
          lut[6916] <= 16'd1211;
          lut[6917] <= 16'd1513;
          lut[6918] <= 16'd1813;
          lut[6919] <= 16'd2112;
          lut[6920] <= 16'd2410;
          lut[6921] <= 16'd2706;
          lut[6922] <= 16'd3000;
          lut[6923] <= 16'd3292;
          lut[6924] <= 16'd3583;
          lut[6925] <= 16'd3871;
          lut[6926] <= 16'd4156;
          lut[6927] <= 16'd4439;
          lut[6928] <= 16'd4720;
          lut[6929] <= 16'd4997;
          lut[6930] <= 16'd5272;
          lut[6931] <= 16'd5543;
          lut[6932] <= 16'd5811;
          lut[6933] <= 16'd6077;
          lut[6934] <= 16'd6339;
          lut[6935] <= 16'd6597;
          lut[6936] <= 16'd6852;
          lut[6937] <= 16'd7104;
          lut[6938] <= 16'd7352;
          lut[6939] <= 16'd7596;
          lut[6940] <= 16'd7837;
          lut[6941] <= 16'd8075;
          lut[6942] <= 16'd8308;
          lut[6943] <= 16'd8538;
          lut[6944] <= 16'd8765;
          lut[6945] <= 16'd8987;
          lut[6946] <= 16'd9207;
          lut[6947] <= 16'd9422;
          lut[6948] <= 16'd9634;
          lut[6949] <= 16'd9842;
          lut[6950] <= 16'd10047;
          lut[6951] <= 16'd10248;
          lut[6952] <= 16'd10446;
          lut[6953] <= 16'd10640;
          lut[6954] <= 16'd10831;
          lut[6955] <= 16'd11018;
          lut[6956] <= 16'd11202;
          lut[6957] <= 16'd11383;
          lut[6958] <= 16'd11560;
          lut[6959] <= 16'd11734;
          lut[6960] <= 16'd11905;
          lut[6961] <= 16'd12073;
          lut[6962] <= 16'd12238;
          lut[6963] <= 16'd12400;
          lut[6964] <= 16'd12559;
          lut[6965] <= 16'd12715;
          lut[6966] <= 16'd12868;
          lut[6967] <= 16'd13018;
          lut[6968] <= 16'd13166;
          lut[6969] <= 16'd13311;
          lut[6970] <= 16'd13453;
          lut[6971] <= 16'd13592;
          lut[6972] <= 16'd13729;
          lut[6973] <= 16'd13864;
          lut[6974] <= 16'd13996;
          lut[6975] <= 16'd14126;
          lut[6976] <= 16'd14253;
          lut[6977] <= 16'd14378;
          lut[6978] <= 16'd14501;
          lut[6979] <= 16'd14622;
          lut[6980] <= 16'd14740;
          lut[6981] <= 16'd14856;
          lut[6982] <= 16'd14970;
          lut[6983] <= 16'd15083;
          lut[6984] <= 16'd15193;
          lut[6985] <= 16'd15301;
          lut[6986] <= 16'd15407;
          lut[6987] <= 16'd15512;
          lut[6988] <= 16'd15615;
          lut[6989] <= 16'd15716;
          lut[6990] <= 16'd15815;
          lut[6991] <= 16'd15912;
          lut[6992] <= 16'd16008;
          lut[6993] <= 16'd16102;
          lut[6994] <= 16'd16195;
          lut[6995] <= 16'd16286;
          lut[6996] <= 16'd16375;
          lut[6997] <= 16'd16463;
          lut[6998] <= 16'd16550;
          lut[6999] <= 16'd16635;
          lut[7000] <= 16'd16718;
          lut[7001] <= 16'd16801;
          lut[7002] <= 16'd16882;
          lut[7003] <= 16'd16961;
          lut[7004] <= 16'd17040;
          lut[7005] <= 16'd17117;
          lut[7006] <= 16'd17193;
          lut[7007] <= 16'd17267;
          lut[7008] <= 16'd17341;
          lut[7009] <= 16'd17413;
          lut[7010] <= 16'd17485;
          lut[7011] <= 16'd17555;
          lut[7012] <= 16'd17624;
          lut[7013] <= 16'd17692;
          lut[7014] <= 16'd17759;
          lut[7015] <= 16'd17824;
          lut[7016] <= 16'd17889;
          lut[7017] <= 16'd17953;
          lut[7018] <= 16'd18016;
          lut[7019] <= 16'd18078;
          lut[7020] <= 16'd18140;
          lut[7021] <= 16'd18200;
          lut[7022] <= 16'd18259;
          lut[7023] <= 16'd18318;
          lut[7024] <= 16'd18375;
          lut[7025] <= 16'd18432;
          lut[7026] <= 16'd18488;
          lut[7027] <= 16'd18543;
          lut[7028] <= 16'd18598;
          lut[7029] <= 16'd18651;
          lut[7030] <= 16'd18704;
          lut[7031] <= 16'd18756;
          lut[7032] <= 16'd18808;
          lut[7033] <= 16'd18859;
          lut[7034] <= 16'd18909;
          lut[7035] <= 16'd18958;
          lut[7036] <= 16'd19007;
          lut[7037] <= 16'd19055;
          lut[7038] <= 16'd19102;
          lut[7039] <= 16'd19149;
          lut[7040] <= 0;
          lut[7041] <= 16'd298;
          lut[7042] <= 16'd596;
          lut[7043] <= 16'd893;
          lut[7044] <= 16'd1189;
          lut[7045] <= 16'd1485;
          lut[7046] <= 16'd1780;
          lut[7047] <= 16'd2074;
          lut[7048] <= 16'd2367;
          lut[7049] <= 16'd2657;
          lut[7050] <= 16'd2947;
          lut[7051] <= 16'd3234;
          lut[7052] <= 16'd3520;
          lut[7053] <= 16'd3803;
          lut[7054] <= 16'd4084;
          lut[7055] <= 16'd4362;
          lut[7056] <= 16'd4638;
          lut[7057] <= 16'd4912;
          lut[7058] <= 16'd5182;
          lut[7059] <= 16'd5450;
          lut[7060] <= 16'd5714;
          lut[7061] <= 16'd5976;
          lut[7062] <= 16'd6234;
          lut[7063] <= 16'd6489;
          lut[7064] <= 16'd6741;
          lut[7065] <= 16'd6990;
          lut[7066] <= 16'd7235;
          lut[7067] <= 16'd7477;
          lut[7068] <= 16'd7715;
          lut[7069] <= 16'd7950;
          lut[7070] <= 16'd8181;
          lut[7071] <= 16'd8409;
          lut[7072] <= 16'd8633;
          lut[7073] <= 16'd8854;
          lut[7074] <= 16'd9072;
          lut[7075] <= 16'd9285;
          lut[7076] <= 16'd9496;
          lut[7077] <= 16'd9702;
          lut[7078] <= 16'd9906;
          lut[7079] <= 16'd10106;
          lut[7080] <= 16'd10302;
          lut[7081] <= 16'd10495;
          lut[7082] <= 16'd10685;
          lut[7083] <= 16'd10872;
          lut[7084] <= 16'd11055;
          lut[7085] <= 16'd11235;
          lut[7086] <= 16'd11412;
          lut[7087] <= 16'd11586;
          lut[7088] <= 16'd11756;
          lut[7089] <= 16'd11924;
          lut[7090] <= 16'd12088;
          lut[7091] <= 16'd12250;
          lut[7092] <= 16'd12409;
          lut[7093] <= 16'd12565;
          lut[7094] <= 16'd12718;
          lut[7095] <= 16'd12868;
          lut[7096] <= 16'd13016;
          lut[7097] <= 16'd13161;
          lut[7098] <= 16'd13303;
          lut[7099] <= 16'd13443;
          lut[7100] <= 16'd13580;
          lut[7101] <= 16'd13715;
          lut[7102] <= 16'd13847;
          lut[7103] <= 16'd13977;
          lut[7104] <= 16'd14105;
          lut[7105] <= 16'd14230;
          lut[7106] <= 16'd14353;
          lut[7107] <= 16'd14474;
          lut[7108] <= 16'd14593;
          lut[7109] <= 16'd14710;
          lut[7110] <= 16'd14825;
          lut[7111] <= 16'd14937;
          lut[7112] <= 16'd15048;
          lut[7113] <= 16'd15157;
          lut[7114] <= 16'd15264;
          lut[7115] <= 16'd15369;
          lut[7116] <= 16'd15472;
          lut[7117] <= 16'd15574;
          lut[7118] <= 16'd15674;
          lut[7119] <= 16'd15772;
          lut[7120] <= 16'd15868;
          lut[7121] <= 16'd15963;
          lut[7122] <= 16'd16056;
          lut[7123] <= 16'd16148;
          lut[7124] <= 16'd16238;
          lut[7125] <= 16'd16327;
          lut[7126] <= 16'd16414;
          lut[7127] <= 16'd16499;
          lut[7128] <= 16'd16584;
          lut[7129] <= 16'd16667;
          lut[7130] <= 16'd16748;
          lut[7131] <= 16'd16829;
          lut[7132] <= 16'd16908;
          lut[7133] <= 16'd16986;
          lut[7134] <= 16'd17062;
          lut[7135] <= 16'd17138;
          lut[7136] <= 16'd17212;
          lut[7137] <= 16'd17285;
          lut[7138] <= 16'd17357;
          lut[7139] <= 16'd17428;
          lut[7140] <= 16'd17497;
          lut[7141] <= 16'd17566;
          lut[7142] <= 16'd17634;
          lut[7143] <= 16'd17700;
          lut[7144] <= 16'd17766;
          lut[7145] <= 16'd17830;
          lut[7146] <= 16'd17894;
          lut[7147] <= 16'd17957;
          lut[7148] <= 16'd18019;
          lut[7149] <= 16'd18080;
          lut[7150] <= 16'd18140;
          lut[7151] <= 16'd18199;
          lut[7152] <= 16'd18257;
          lut[7153] <= 16'd18314;
          lut[7154] <= 16'd18371;
          lut[7155] <= 16'd18427;
          lut[7156] <= 16'd18482;
          lut[7157] <= 16'd18536;
          lut[7158] <= 16'd18590;
          lut[7159] <= 16'd18643;
          lut[7160] <= 16'd18695;
          lut[7161] <= 16'd18746;
          lut[7162] <= 16'd18797;
          lut[7163] <= 16'd18847;
          lut[7164] <= 16'd18896;
          lut[7165] <= 16'd18945;
          lut[7166] <= 16'd18993;
          lut[7167] <= 16'd19040;
          lut[7168] <= 0;
          lut[7169] <= 16'd293;
          lut[7170] <= 16'd585;
          lut[7171] <= 16'd877;
          lut[7172] <= 16'd1168;
          lut[7173] <= 16'd1459;
          lut[7174] <= 16'd1749;
          lut[7175] <= 16'd2037;
          lut[7176] <= 16'd2325;
          lut[7177] <= 16'd2611;
          lut[7178] <= 16'd2895;
          lut[7179] <= 16'd3178;
          lut[7180] <= 16'd3459;
          lut[7181] <= 16'd3737;
          lut[7182] <= 16'd4014;
          lut[7183] <= 16'd4288;
          lut[7184] <= 16'd4560;
          lut[7185] <= 16'd4829;
          lut[7186] <= 16'd5095;
          lut[7187] <= 16'd5359;
          lut[7188] <= 16'd5620;
          lut[7189] <= 16'd5878;
          lut[7190] <= 16'd6133;
          lut[7191] <= 16'd6385;
          lut[7192] <= 16'd6634;
          lut[7193] <= 16'd6879;
          lut[7194] <= 16'd7122;
          lut[7195] <= 16'd7361;
          lut[7196] <= 16'd7596;
          lut[7197] <= 16'd7829;
          lut[7198] <= 16'd8058;
          lut[7199] <= 16'd8283;
          lut[7200] <= 16'd8506;
          lut[7201] <= 16'd8725;
          lut[7202] <= 16'd8940;
          lut[7203] <= 16'd9152;
          lut[7204] <= 16'd9361;
          lut[7205] <= 16'd9566;
          lut[7206] <= 16'd9768;
          lut[7207] <= 16'd9967;
          lut[7208] <= 16'd10162;
          lut[7209] <= 16'd10354;
          lut[7210] <= 16'd10543;
          lut[7211] <= 16'd10729;
          lut[7212] <= 16'd10911;
          lut[7213] <= 16'd11091;
          lut[7214] <= 16'd11267;
          lut[7215] <= 16'd11440;
          lut[7216] <= 16'd11610;
          lut[7217] <= 16'd11777;
          lut[7218] <= 16'd11942;
          lut[7219] <= 16'd12103;
          lut[7220] <= 16'd12261;
          lut[7221] <= 16'd12417;
          lut[7222] <= 16'd12570;
          lut[7223] <= 16'd12720;
          lut[7224] <= 16'd12868;
          lut[7225] <= 16'd13013;
          lut[7226] <= 16'd13155;
          lut[7227] <= 16'd13295;
          lut[7228] <= 16'd13433;
          lut[7229] <= 16'd13568;
          lut[7230] <= 16'd13700;
          lut[7231] <= 16'd13831;
          lut[7232] <= 16'd13959;
          lut[7233] <= 16'd14084;
          lut[7234] <= 16'd14208;
          lut[7235] <= 16'd14329;
          lut[7236] <= 16'd14449;
          lut[7237] <= 16'd14566;
          lut[7238] <= 16'd14681;
          lut[7239] <= 16'd14794;
          lut[7240] <= 16'd14905;
          lut[7241] <= 16'd15015;
          lut[7242] <= 16'd15122;
          lut[7243] <= 16'd15228;
          lut[7244] <= 16'd15332;
          lut[7245] <= 16'd15434;
          lut[7246] <= 16'd15534;
          lut[7247] <= 16'd15633;
          lut[7248] <= 16'd15730;
          lut[7249] <= 16'd15825;
          lut[7250] <= 16'd15919;
          lut[7251] <= 16'd16011;
          lut[7252] <= 16'd16102;
          lut[7253] <= 16'd16191;
          lut[7254] <= 16'd16279;
          lut[7255] <= 16'd16366;
          lut[7256] <= 16'd16451;
          lut[7257] <= 16'd16534;
          lut[7258] <= 16'd16617;
          lut[7259] <= 16'd16698;
          lut[7260] <= 16'd16777;
          lut[7261] <= 16'd16856;
          lut[7262] <= 16'd16933;
          lut[7263] <= 16'd17009;
          lut[7264] <= 16'd17084;
          lut[7265] <= 16'd17158;
          lut[7266] <= 16'd17230;
          lut[7267] <= 16'd17302;
          lut[7268] <= 16'd17372;
          lut[7269] <= 16'd17441;
          lut[7270] <= 16'd17510;
          lut[7271] <= 16'd17577;
          lut[7272] <= 16'd17643;
          lut[7273] <= 16'd17708;
          lut[7274] <= 16'd17773;
          lut[7275] <= 16'd17836;
          lut[7276] <= 16'd17899;
          lut[7277] <= 16'd17960;
          lut[7278] <= 16'd18021;
          lut[7279] <= 16'd18081;
          lut[7280] <= 16'd18140;
          lut[7281] <= 16'd18198;
          lut[7282] <= 16'd18255;
          lut[7283] <= 16'd18311;
          lut[7284] <= 16'd18367;
          lut[7285] <= 16'd18422;
          lut[7286] <= 16'd18476;
          lut[7287] <= 16'd18530;
          lut[7288] <= 16'd18582;
          lut[7289] <= 16'd18634;
          lut[7290] <= 16'd18685;
          lut[7291] <= 16'd18736;
          lut[7292] <= 16'd18786;
          lut[7293] <= 16'd18835;
          lut[7294] <= 16'd18884;
          lut[7295] <= 16'd18932;
          lut[7296] <= 0;
          lut[7297] <= 16'd287;
          lut[7298] <= 16'd575;
          lut[7299] <= 16'd862;
          lut[7300] <= 16'd1148;
          lut[7301] <= 16'd1434;
          lut[7302] <= 16'd1718;
          lut[7303] <= 16'd2002;
          lut[7304] <= 16'd2285;
          lut[7305] <= 16'd2566;
          lut[7306] <= 16'd2845;
          lut[7307] <= 16'd3123;
          lut[7308] <= 16'd3400;
          lut[7309] <= 16'd3674;
          lut[7310] <= 16'd3946;
          lut[7311] <= 16'd4216;
          lut[7312] <= 16'd4484;
          lut[7313] <= 16'd4749;
          lut[7314] <= 16'd5012;
          lut[7315] <= 16'd5272;
          lut[7316] <= 16'd5529;
          lut[7317] <= 16'd5783;
          lut[7318] <= 16'd6035;
          lut[7319] <= 16'd6284;
          lut[7320] <= 16'd6529;
          lut[7321] <= 16'd6772;
          lut[7322] <= 16'd7012;
          lut[7323] <= 16'd7248;
          lut[7324] <= 16'd7481;
          lut[7325] <= 16'd7711;
          lut[7326] <= 16'd7938;
          lut[7327] <= 16'd8161;
          lut[7328] <= 16'd8381;
          lut[7329] <= 16'd8598;
          lut[7330] <= 16'd8812;
          lut[7331] <= 16'd9022;
          lut[7332] <= 16'd9229;
          lut[7333] <= 16'd9433;
          lut[7334] <= 16'd9634;
          lut[7335] <= 16'd9831;
          lut[7336] <= 16'd10025;
          lut[7337] <= 16'd10216;
          lut[7338] <= 16'd10404;
          lut[7339] <= 16'd10589;
          lut[7340] <= 16'd10771;
          lut[7341] <= 16'd10949;
          lut[7342] <= 16'd11125;
          lut[7343] <= 16'd11297;
          lut[7344] <= 16'd11467;
          lut[7345] <= 16'd11634;
          lut[7346] <= 16'd11798;
          lut[7347] <= 16'd11959;
          lut[7348] <= 16'd12117;
          lut[7349] <= 16'd12272;
          lut[7350] <= 16'd12425;
          lut[7351] <= 16'd12575;
          lut[7352] <= 16'd12723;
          lut[7353] <= 16'd12868;
          lut[7354] <= 16'd13010;
          lut[7355] <= 16'd13150;
          lut[7356] <= 16'd13288;
          lut[7357] <= 16'd13423;
          lut[7358] <= 16'd13556;
          lut[7359] <= 16'd13686;
          lut[7360] <= 16'd13815;
          lut[7361] <= 16'd13941;
          lut[7362] <= 16'd14065;
          lut[7363] <= 16'd14186;
          lut[7364] <= 16'd14306;
          lut[7365] <= 16'd14424;
          lut[7366] <= 16'd14539;
          lut[7367] <= 16'd14653;
          lut[7368] <= 16'd14765;
          lut[7369] <= 16'd14874;
          lut[7370] <= 16'd14982;
          lut[7371] <= 16'd15088;
          lut[7372] <= 16'd15193;
          lut[7373] <= 16'd15295;
          lut[7374] <= 16'd15396;
          lut[7375] <= 16'd15496;
          lut[7376] <= 16'd15593;
          lut[7377] <= 16'd15689;
          lut[7378] <= 16'd15784;
          lut[7379] <= 16'd15876;
          lut[7380] <= 16'd15968;
          lut[7381] <= 16'd16058;
          lut[7382] <= 16'd16146;
          lut[7383] <= 16'd16233;
          lut[7384] <= 16'd16319;
          lut[7385] <= 16'd16403;
          lut[7386] <= 16'd16486;
          lut[7387] <= 16'd16568;
          lut[7388] <= 16'd16648;
          lut[7389] <= 16'd16727;
          lut[7390] <= 16'd16805;
          lut[7391] <= 16'd16882;
          lut[7392] <= 16'd16957;
          lut[7393] <= 16'd17032;
          lut[7394] <= 16'd17105;
          lut[7395] <= 16'd17177;
          lut[7396] <= 16'd17248;
          lut[7397] <= 16'd17318;
          lut[7398] <= 16'd17387;
          lut[7399] <= 16'd17455;
          lut[7400] <= 16'd17522;
          lut[7401] <= 16'd17587;
          lut[7402] <= 16'd17652;
          lut[7403] <= 16'd17716;
          lut[7404] <= 16'd17779;
          lut[7405] <= 16'd17842;
          lut[7406] <= 16'd17903;
          lut[7407] <= 16'd17963;
          lut[7408] <= 16'd18023;
          lut[7409] <= 16'd18082;
          lut[7410] <= 16'd18140;
          lut[7411] <= 16'd18197;
          lut[7412] <= 16'd18253;
          lut[7413] <= 16'd18308;
          lut[7414] <= 16'd18363;
          lut[7415] <= 16'd18417;
          lut[7416] <= 16'd18470;
          lut[7417] <= 16'd18523;
          lut[7418] <= 16'd18575;
          lut[7419] <= 16'd18626;
          lut[7420] <= 16'd18677;
          lut[7421] <= 16'd18726;
          lut[7422] <= 16'd18775;
          lut[7423] <= 16'd18824;
          lut[7424] <= 0;
          lut[7425] <= 16'd282;
          lut[7426] <= 16'd565;
          lut[7427] <= 16'd847;
          lut[7428] <= 16'd1128;
          lut[7429] <= 16'd1409;
          lut[7430] <= 16'd1689;
          lut[7431] <= 16'd1968;
          lut[7432] <= 16'd2246;
          lut[7433] <= 16'd2522;
          lut[7434] <= 16'd2797;
          lut[7435] <= 16'd3071;
          lut[7436] <= 16'd3343;
          lut[7437] <= 16'd3613;
          lut[7438] <= 16'd3881;
          lut[7439] <= 16'd4146;
          lut[7440] <= 16'd4410;
          lut[7441] <= 16'd4671;
          lut[7442] <= 16'd4930;
          lut[7443] <= 16'd5187;
          lut[7444] <= 16'd5440;
          lut[7445] <= 16'd5692;
          lut[7446] <= 16'd5940;
          lut[7447] <= 16'd6185;
          lut[7448] <= 16'd6428;
          lut[7449] <= 16'd6668;
          lut[7450] <= 16'd6905;
          lut[7451] <= 16'd7138;
          lut[7452] <= 16'd7369;
          lut[7453] <= 16'd7596;
          lut[7454] <= 16'd7821;
          lut[7455] <= 16'd8042;
          lut[7456] <= 16'd8260;
          lut[7457] <= 16'd8475;
          lut[7458] <= 16'd8687;
          lut[7459] <= 16'd8896;
          lut[7460] <= 16'd9101;
          lut[7461] <= 16'd9304;
          lut[7462] <= 16'd9503;
          lut[7463] <= 16'd9699;
          lut[7464] <= 16'd9892;
          lut[7465] <= 16'd10082;
          lut[7466] <= 16'd10269;
          lut[7467] <= 16'd10452;
          lut[7468] <= 16'd10633;
          lut[7469] <= 16'd10811;
          lut[7470] <= 16'd10986;
          lut[7471] <= 16'd11158;
          lut[7472] <= 16'd11327;
          lut[7473] <= 16'd11493;
          lut[7474] <= 16'd11657;
          lut[7475] <= 16'd11817;
          lut[7476] <= 16'd11975;
          lut[7477] <= 16'd12130;
          lut[7478] <= 16'd12283;
          lut[7479] <= 16'd12433;
          lut[7480] <= 16'd12581;
          lut[7481] <= 16'd12725;
          lut[7482] <= 16'd12868;
          lut[7483] <= 16'd13008;
          lut[7484] <= 16'd13146;
          lut[7485] <= 16'd13281;
          lut[7486] <= 16'd13414;
          lut[7487] <= 16'd13545;
          lut[7488] <= 16'd13673;
          lut[7489] <= 16'd13799;
          lut[7490] <= 16'd13924;
          lut[7491] <= 16'd14046;
          lut[7492] <= 16'd14166;
          lut[7493] <= 16'd14284;
          lut[7494] <= 16'd14399;
          lut[7495] <= 16'd14514;
          lut[7496] <= 16'd14626;
          lut[7497] <= 16'd14736;
          lut[7498] <= 16'd14844;
          lut[7499] <= 16'd14951;
          lut[7500] <= 16'd15056;
          lut[7501] <= 16'd15159;
          lut[7502] <= 16'd15260;
          lut[7503] <= 16'd15360;
          lut[7504] <= 16'd15458;
          lut[7505] <= 16'd15555;
          lut[7506] <= 16'd15650;
          lut[7507] <= 16'd15743;
          lut[7508] <= 16'd15835;
          lut[7509] <= 16'd15925;
          lut[7510] <= 16'd16014;
          lut[7511] <= 16'd16102;
          lut[7512] <= 16'd16188;
          lut[7513] <= 16'd16273;
          lut[7514] <= 16'd16357;
          lut[7515] <= 16'd16439;
          lut[7516] <= 16'd16520;
          lut[7517] <= 16'd16600;
          lut[7518] <= 16'd16678;
          lut[7519] <= 16'd16755;
          lut[7520] <= 16'd16832;
          lut[7521] <= 16'd16907;
          lut[7522] <= 16'd16980;
          lut[7523] <= 16'd17053;
          lut[7524] <= 16'd17125;
          lut[7525] <= 16'd17195;
          lut[7526] <= 16'd17265;
          lut[7527] <= 16'd17333;
          lut[7528] <= 16'd17401;
          lut[7529] <= 16'd17467;
          lut[7530] <= 16'd17533;
          lut[7531] <= 16'd17598;
          lut[7532] <= 16'd17661;
          lut[7533] <= 16'd17724;
          lut[7534] <= 16'd17786;
          lut[7535] <= 16'd17847;
          lut[7536] <= 16'd17907;
          lut[7537] <= 16'd17966;
          lut[7538] <= 16'd18025;
          lut[7539] <= 16'd18083;
          lut[7540] <= 16'd18140;
          lut[7541] <= 16'd18196;
          lut[7542] <= 16'd18251;
          lut[7543] <= 16'd18306;
          lut[7544] <= 16'd18359;
          lut[7545] <= 16'd18413;
          lut[7546] <= 16'd18465;
          lut[7547] <= 16'd18517;
          lut[7548] <= 16'd18568;
          lut[7549] <= 16'd18618;
          lut[7550] <= 16'd18668;
          lut[7551] <= 16'd18717;
          lut[7552] <= 0;
          lut[7553] <= 16'd278;
          lut[7554] <= 16'd555;
          lut[7555] <= 16'd832;
          lut[7556] <= 16'd1109;
          lut[7557] <= 16'd1385;
          lut[7558] <= 16'd1660;
          lut[7559] <= 16'd1935;
          lut[7560] <= 16'd2208;
          lut[7561] <= 16'd2480;
          lut[7562] <= 16'd2751;
          lut[7563] <= 16'd3020;
          lut[7564] <= 16'd3287;
          lut[7565] <= 16'd3553;
          lut[7566] <= 16'd3817;
          lut[7567] <= 16'd4079;
          lut[7568] <= 16'd4339;
          lut[7569] <= 16'd4596;
          lut[7570] <= 16'd4852;
          lut[7571] <= 16'd5104;
          lut[7572] <= 16'd5355;
          lut[7573] <= 16'd5603;
          lut[7574] <= 16'd5848;
          lut[7575] <= 16'd6090;
          lut[7576] <= 16'd6330;
          lut[7577] <= 16'd6567;
          lut[7578] <= 16'd6801;
          lut[7579] <= 16'd7032;
          lut[7580] <= 16'd7260;
          lut[7581] <= 16'd7485;
          lut[7582] <= 16'd7707;
          lut[7583] <= 16'd7926;
          lut[7584] <= 16'd8142;
          lut[7585] <= 16'd8355;
          lut[7586] <= 16'd8565;
          lut[7587] <= 16'd8772;
          lut[7588] <= 16'd8976;
          lut[7589] <= 16'd9177;
          lut[7590] <= 16'd9375;
          lut[7591] <= 16'd9570;
          lut[7592] <= 16'd9761;
          lut[7593] <= 16'd9950;
          lut[7594] <= 16'd10136;
          lut[7595] <= 16'd10319;
          lut[7596] <= 16'd10499;
          lut[7597] <= 16'd10676;
          lut[7598] <= 16'd10850;
          lut[7599] <= 16'd11021;
          lut[7600] <= 16'd11190;
          lut[7601] <= 16'd11355;
          lut[7602] <= 16'd11518;
          lut[7603] <= 16'd11678;
          lut[7604] <= 16'd11836;
          lut[7605] <= 16'd11991;
          lut[7606] <= 16'd12143;
          lut[7607] <= 16'd12293;
          lut[7608] <= 16'd12441;
          lut[7609] <= 16'd12586;
          lut[7610] <= 16'd12728;
          lut[7611] <= 16'd12868;
          lut[7612] <= 16'd13006;
          lut[7613] <= 16'd13141;
          lut[7614] <= 16'd13274;
          lut[7615] <= 16'd13405;
          lut[7616] <= 16'd13534;
          lut[7617] <= 16'd13660;
          lut[7618] <= 16'd13785;
          lut[7619] <= 16'd13907;
          lut[7620] <= 16'd14027;
          lut[7621] <= 16'd14145;
          lut[7622] <= 16'd14262;
          lut[7623] <= 16'd14376;
          lut[7624] <= 16'd14489;
          lut[7625] <= 16'd14599;
          lut[7626] <= 16'd14708;
          lut[7627] <= 16'd14815;
          lut[7628] <= 16'd14920;
          lut[7629] <= 16'd15024;
          lut[7630] <= 16'd15126;
          lut[7631] <= 16'd15226;
          lut[7632] <= 16'd15325;
          lut[7633] <= 16'd15422;
          lut[7634] <= 16'd15517;
          lut[7635] <= 16'd15611;
          lut[7636] <= 16'd15704;
          lut[7637] <= 16'd15795;
          lut[7638] <= 16'd15884;
          lut[7639] <= 16'd15972;
          lut[7640] <= 16'd16059;
          lut[7641] <= 16'd16145;
          lut[7642] <= 16'd16229;
          lut[7643] <= 16'd16312;
          lut[7644] <= 16'd16393;
          lut[7645] <= 16'd16473;
          lut[7646] <= 16'd16553;
          lut[7647] <= 16'd16630;
          lut[7648] <= 16'd16707;
          lut[7649] <= 16'd16783;
          lut[7650] <= 16'd16857;
          lut[7651] <= 16'd16930;
          lut[7652] <= 16'd17003;
          lut[7653] <= 16'd17074;
          lut[7654] <= 16'd17144;
          lut[7655] <= 16'd17213;
          lut[7656] <= 16'd17281;
          lut[7657] <= 16'd17348;
          lut[7658] <= 16'd17415;
          lut[7659] <= 16'd17480;
          lut[7660] <= 16'd17544;
          lut[7661] <= 16'd17607;
          lut[7662] <= 16'd17670;
          lut[7663] <= 16'd17731;
          lut[7664] <= 16'd17792;
          lut[7665] <= 16'd17852;
          lut[7666] <= 16'd17911;
          lut[7667] <= 16'd17969;
          lut[7668] <= 16'd18027;
          lut[7669] <= 16'd18084;
          lut[7670] <= 16'd18140;
          lut[7671] <= 16'd18195;
          lut[7672] <= 16'd18249;
          lut[7673] <= 16'd18303;
          lut[7674] <= 16'd18356;
          lut[7675] <= 16'd18408;
          lut[7676] <= 16'd18460;
          lut[7677] <= 16'd18511;
          lut[7678] <= 16'd18561;
          lut[7679] <= 16'd18611;
          lut[7680] <= 0;
          lut[7681] <= 16'd273;
          lut[7682] <= 16'd546;
          lut[7683] <= 16'd819;
          lut[7684] <= 16'd1091;
          lut[7685] <= 16'd1362;
          lut[7686] <= 16'd1633;
          lut[7687] <= 16'd1903;
          lut[7688] <= 16'd2172;
          lut[7689] <= 16'd2439;
          lut[7690] <= 16'd2706;
          lut[7691] <= 16'd2971;
          lut[7692] <= 16'd3234;
          lut[7693] <= 16'd3496;
          lut[7694] <= 16'd3756;
          lut[7695] <= 16'd4014;
          lut[7696] <= 16'd4270;
          lut[7697] <= 16'd4524;
          lut[7698] <= 16'd4775;
          lut[7699] <= 16'd5025;
          lut[7700] <= 16'd5272;
          lut[7701] <= 16'd5516;
          lut[7702] <= 16'd5758;
          lut[7703] <= 16'd5997;
          lut[7704] <= 16'd6234;
          lut[7705] <= 16'd6468;
          lut[7706] <= 16'd6700;
          lut[7707] <= 16'd6928;
          lut[7708] <= 16'd7154;
          lut[7709] <= 16'd7376;
          lut[7710] <= 16'd7596;
          lut[7711] <= 16'd7813;
          lut[7712] <= 16'd8027;
          lut[7713] <= 16'd8239;
          lut[7714] <= 16'd8447;
          lut[7715] <= 16'd8652;
          lut[7716] <= 16'd8854;
          lut[7717] <= 16'd9054;
          lut[7718] <= 16'd9250;
          lut[7719] <= 16'd9443;
          lut[7720] <= 16'd9634;
          lut[7721] <= 16'd9821;
          lut[7722] <= 16'd10006;
          lut[7723] <= 16'd10188;
          lut[7724] <= 16'd10367;
          lut[7725] <= 16'd10543;
          lut[7726] <= 16'd10716;
          lut[7727] <= 16'd10887;
          lut[7728] <= 16'd11055;
          lut[7729] <= 16'd11220;
          lut[7730] <= 16'd11383;
          lut[7731] <= 16'd11542;
          lut[7732] <= 16'd11700;
          lut[7733] <= 16'd11854;
          lut[7734] <= 16'd12006;
          lut[7735] <= 16'd12156;
          lut[7736] <= 16'd12303;
          lut[7737] <= 16'd12448;
          lut[7738] <= 16'd12590;
          lut[7739] <= 16'd12730;
          lut[7740] <= 16'd12868;
          lut[7741] <= 16'd13003;
          lut[7742] <= 16'd13137;
          lut[7743] <= 16'd13267;
          lut[7744] <= 16'd13396;
          lut[7745] <= 16'd13523;
          lut[7746] <= 16'd13648;
          lut[7747] <= 16'd13770;
          lut[7748] <= 16'd13891;
          lut[7749] <= 16'd14009;
          lut[7750] <= 16'd14126;
          lut[7751] <= 16'd14240;
          lut[7752] <= 16'd14353;
          lut[7753] <= 16'd14464;
          lut[7754] <= 16'd14574;
          lut[7755] <= 16'd14681;
          lut[7756] <= 16'd14787;
          lut[7757] <= 16'd14891;
          lut[7758] <= 16'd14993;
          lut[7759] <= 16'd15094;
          lut[7760] <= 16'd15193;
          lut[7761] <= 16'd15290;
          lut[7762] <= 16'd15386;
          lut[7763] <= 16'd15481;
          lut[7764] <= 16'd15574;
          lut[7765] <= 16'd15665;
          lut[7766] <= 16'd15755;
          lut[7767] <= 16'd15844;
          lut[7768] <= 16'd15931;
          lut[7769] <= 16'd16017;
          lut[7770] <= 16'd16102;
          lut[7771] <= 16'd16185;
          lut[7772] <= 16'd16268;
          lut[7773] <= 16'd16348;
          lut[7774] <= 16'd16428;
          lut[7775] <= 16'd16507;
          lut[7776] <= 16'd16584;
          lut[7777] <= 16'd16660;
          lut[7778] <= 16'd16735;
          lut[7779] <= 16'd16809;
          lut[7780] <= 16'd16882;
          lut[7781] <= 16'd16953;
          lut[7782] <= 16'd17024;
          lut[7783] <= 16'd17094;
          lut[7784] <= 16'd17163;
          lut[7785] <= 16'd17230;
          lut[7786] <= 16'd17297;
          lut[7787] <= 16'd17363;
          lut[7788] <= 16'd17428;
          lut[7789] <= 16'd17492;
          lut[7790] <= 16'd17555;
          lut[7791] <= 16'd17617;
          lut[7792] <= 16'd17678;
          lut[7793] <= 16'd17739;
          lut[7794] <= 16'd17798;
          lut[7795] <= 16'd17857;
          lut[7796] <= 16'd17915;
          lut[7797] <= 16'd17972;
          lut[7798] <= 16'd18029;
          lut[7799] <= 16'd18085;
          lut[7800] <= 16'd18140;
          lut[7801] <= 16'd18194;
          lut[7802] <= 16'd18247;
          lut[7803] <= 16'd18300;
          lut[7804] <= 16'd18352;
          lut[7805] <= 16'd18404;
          lut[7806] <= 16'd18455;
          lut[7807] <= 16'd18505;
          lut[7808] <= 0;
          lut[7809] <= 16'd269;
          lut[7810] <= 16'd537;
          lut[7811] <= 16'd805;
          lut[7812] <= 16'd1073;
          lut[7813] <= 16'd1340;
          lut[7814] <= 16'd1606;
          lut[7815] <= 16'd1872;
          lut[7816] <= 16'd2137;
          lut[7817] <= 16'd2400;
          lut[7818] <= 16'd2662;
          lut[7819] <= 16'd2923;
          lut[7820] <= 16'd3182;
          lut[7821] <= 16'd3440;
          lut[7822] <= 16'd3696;
          lut[7823] <= 16'd3950;
          lut[7824] <= 16'd4203;
          lut[7825] <= 16'd4453;
          lut[7826] <= 16'd4701;
          lut[7827] <= 16'd4947;
          lut[7828] <= 16'd5191;
          lut[7829] <= 16'd5432;
          lut[7830] <= 16'd5671;
          lut[7831] <= 16'd5908;
          lut[7832] <= 16'd6141;
          lut[7833] <= 16'd6373;
          lut[7834] <= 16'd6601;
          lut[7835] <= 16'd6827;
          lut[7836] <= 16'd7050;
          lut[7837] <= 16'd7271;
          lut[7838] <= 16'd7489;
          lut[7839] <= 16'd7703;
          lut[7840] <= 16'd7916;
          lut[7841] <= 16'd8125;
          lut[7842] <= 16'd8331;
          lut[7843] <= 16'd8535;
          lut[7844] <= 16'd8735;
          lut[7845] <= 16'd8933;
          lut[7846] <= 16'd9128;
          lut[7847] <= 16'd9320;
          lut[7848] <= 16'd9509;
          lut[7849] <= 16'd9696;
          lut[7850] <= 16'd9879;
          lut[7851] <= 16'd10060;
          lut[7852] <= 16'd10238;
          lut[7853] <= 16'd10413;
          lut[7854] <= 16'd10586;
          lut[7855] <= 16'd10756;
          lut[7856] <= 16'd10923;
          lut[7857] <= 16'd11088;
          lut[7858] <= 16'd11250;
          lut[7859] <= 16'd11409;
          lut[7860] <= 16'd11566;
          lut[7861] <= 16'd11720;
          lut[7862] <= 16'd11872;
          lut[7863] <= 16'd12021;
          lut[7864] <= 16'd12168;
          lut[7865] <= 16'd12313;
          lut[7866] <= 16'd12455;
          lut[7867] <= 16'd12595;
          lut[7868] <= 16'd12733;
          lut[7869] <= 16'd12868;
          lut[7870] <= 16'd13001;
          lut[7871] <= 16'd13132;
          lut[7872] <= 16'd13261;
          lut[7873] <= 16'd13388;
          lut[7874] <= 16'd13513;
          lut[7875] <= 16'd13635;
          lut[7876] <= 16'd13756;
          lut[7877] <= 16'd13875;
          lut[7878] <= 16'd13992;
          lut[7879] <= 16'd14107;
          lut[7880] <= 16'd14220;
          lut[7881] <= 16'd14331;
          lut[7882] <= 16'd14441;
          lut[7883] <= 16'd14549;
          lut[7884] <= 16'd14655;
          lut[7885] <= 16'd14759;
          lut[7886] <= 16'd14862;
          lut[7887] <= 16'd14963;
          lut[7888] <= 16'd15063;
          lut[7889] <= 16'd15160;
          lut[7890] <= 16'd15257;
          lut[7891] <= 16'd15352;
          lut[7892] <= 16'd15445;
          lut[7893] <= 16'd15537;
          lut[7894] <= 16'd15628;
          lut[7895] <= 16'd15717;
          lut[7896] <= 16'd15805;
          lut[7897] <= 16'd15892;
          lut[7898] <= 16'd15977;
          lut[7899] <= 16'd16061;
          lut[7900] <= 16'd16143;
          lut[7901] <= 16'd16225;
          lut[7902] <= 16'd16305;
          lut[7903] <= 16'd16384;
          lut[7904] <= 16'd16462;
          lut[7905] <= 16'd16538;
          lut[7906] <= 16'd16614;
          lut[7907] <= 16'd16688;
          lut[7908] <= 16'd16762;
          lut[7909] <= 16'd16834;
          lut[7910] <= 16'd16905;
          lut[7911] <= 16'd16976;
          lut[7912] <= 16'd17045;
          lut[7913] <= 16'd17113;
          lut[7914] <= 16'd17180;
          lut[7915] <= 16'd17247;
          lut[7916] <= 16'd17312;
          lut[7917] <= 16'd17377;
          lut[7918] <= 16'd17440;
          lut[7919] <= 16'd17503;
          lut[7920] <= 16'd17565;
          lut[7921] <= 16'd17626;
          lut[7922] <= 16'd17686;
          lut[7923] <= 16'd17745;
          lut[7924] <= 16'd17804;
          lut[7925] <= 16'd17862;
          lut[7926] <= 16'd17919;
          lut[7927] <= 16'd17975;
          lut[7928] <= 16'd18031;
          lut[7929] <= 16'd18085;
          lut[7930] <= 16'd18140;
          lut[7931] <= 16'd18193;
          lut[7932] <= 16'd18246;
          lut[7933] <= 16'd18298;
          lut[7934] <= 16'd18349;
          lut[7935] <= 16'd18400;
          lut[7936] <= 0;
          lut[7937] <= 16'd264;
          lut[7938] <= 16'd528;
          lut[7939] <= 16'd792;
          lut[7940] <= 16'd1056;
          lut[7941] <= 16'd1318;
          lut[7942] <= 16'd1581;
          lut[7943] <= 16'd1842;
          lut[7944] <= 16'd2102;
          lut[7945] <= 16'd2362;
          lut[7946] <= 16'd2620;
          lut[7947] <= 16'd2877;
          lut[7948] <= 16'd3132;
          lut[7949] <= 16'd3386;
          lut[7950] <= 16'd3639;
          lut[7951] <= 16'd3889;
          lut[7952] <= 16'd4138;
          lut[7953] <= 16'd4385;
          lut[7954] <= 16'd4629;
          lut[7955] <= 16'd4872;
          lut[7956] <= 16'd5112;
          lut[7957] <= 16'd5351;
          lut[7958] <= 16'd5587;
          lut[7959] <= 16'd5820;
          lut[7960] <= 16'd6051;
          lut[7961] <= 16'd6280;
          lut[7962] <= 16'd6506;
          lut[7963] <= 16'd6729;
          lut[7964] <= 16'd6950;
          lut[7965] <= 16'd7168;
          lut[7966] <= 16'd7384;
          lut[7967] <= 16'd7596;
          lut[7968] <= 16'd7806;
          lut[7969] <= 16'd8014;
          lut[7970] <= 16'd8218;
          lut[7971] <= 16'd8420;
          lut[7972] <= 16'd8619;
          lut[7973] <= 16'd8815;
          lut[7974] <= 16'd9009;
          lut[7975] <= 16'd9200;
          lut[7976] <= 16'd9387;
          lut[7977] <= 16'd9573;
          lut[7978] <= 16'd9755;
          lut[7979] <= 16'd9935;
          lut[7980] <= 16'd10112;
          lut[7981] <= 16'd10286;
          lut[7982] <= 16'd10458;
          lut[7983] <= 16'd10627;
          lut[7984] <= 16'd10794;
          lut[7985] <= 16'd10958;
          lut[7986] <= 16'd11119;
          lut[7987] <= 16'd11278;
          lut[7988] <= 16'd11434;
          lut[7989] <= 16'd11588;
          lut[7990] <= 16'd11740;
          lut[7991] <= 16'd11889;
          lut[7992] <= 16'd12036;
          lut[7993] <= 16'd12180;
          lut[7994] <= 16'd12322;
          lut[7995] <= 16'd12462;
          lut[7996] <= 16'd12599;
          lut[7997] <= 16'd12735;
          lut[7998] <= 16'd12868;
          lut[7999] <= 16'd12999;
          lut[8000] <= 16'd13128;
          lut[8001] <= 16'd13255;
          lut[8002] <= 16'd13380;
          lut[8003] <= 16'd13503;
          lut[8004] <= 16'd13624;
          lut[8005] <= 16'd13743;
          lut[8006] <= 16'd13860;
          lut[8007] <= 16'd13975;
          lut[8008] <= 16'd14088;
          lut[8009] <= 16'd14200;
          lut[8010] <= 16'd14310;
          lut[8011] <= 16'd14418;
          lut[8012] <= 16'd14524;
          lut[8013] <= 16'd14629;
          lut[8014] <= 16'd14732;
          lut[8015] <= 16'd14834;
          lut[8016] <= 16'd14934;
          lut[8017] <= 16'd15032;
          lut[8018] <= 16'd15129;
          lut[8019] <= 16'd15224;
          lut[8020] <= 16'd15318;
          lut[8021] <= 16'd15411;
          lut[8022] <= 16'd15502;
          lut[8023] <= 16'd15592;
          lut[8024] <= 16'd15680;
          lut[8025] <= 16'd15767;
          lut[8026] <= 16'd15853;
          lut[8027] <= 16'd15937;
          lut[8028] <= 16'd16020;
          lut[8029] <= 16'd16102;
          lut[8030] <= 16'd16183;
          lut[8031] <= 16'd16262;
          lut[8032] <= 16'd16341;
          lut[8033] <= 16'd16418;
          lut[8034] <= 16'd16494;
          lut[8035] <= 16'd16569;
          lut[8036] <= 16'd16643;
          lut[8037] <= 16'd16716;
          lut[8038] <= 16'd16788;
          lut[8039] <= 16'd16858;
          lut[8040] <= 16'd16928;
          lut[8041] <= 16'd16997;
          lut[8042] <= 16'd17065;
          lut[8043] <= 16'd17132;
          lut[8044] <= 16'd17198;
          lut[8045] <= 16'd17263;
          lut[8046] <= 16'd17327;
          lut[8047] <= 16'd17390;
          lut[8048] <= 16'd17452;
          lut[8049] <= 16'd17514;
          lut[8050] <= 16'd17575;
          lut[8051] <= 16'd17635;
          lut[8052] <= 16'd17694;
          lut[8053] <= 16'd17752;
          lut[8054] <= 16'd17810;
          lut[8055] <= 16'd17866;
          lut[8056] <= 16'd17923;
          lut[8057] <= 16'd17978;
          lut[8058] <= 16'd18032;
          lut[8059] <= 16'd18086;
          lut[8060] <= 16'd18140;
          lut[8061] <= 16'd18192;
          lut[8062] <= 16'd18244;
          lut[8063] <= 16'd18295;
          lut[8064] <= 0;
          lut[8065] <= 16'd260;
          lut[8066] <= 16'd520;
          lut[8067] <= 16'd780;
          lut[8068] <= 16'd1039;
          lut[8069] <= 16'd1298;
          lut[8070] <= 16'd1556;
          lut[8071] <= 16'd1813;
          lut[8072] <= 16'd2069;
          lut[8073] <= 16'd2325;
          lut[8074] <= 16'd2579;
          lut[8075] <= 16'd2832;
          lut[8076] <= 16'd3084;
          lut[8077] <= 16'd3334;
          lut[8078] <= 16'd3583;
          lut[8079] <= 16'd3830;
          lut[8080] <= 16'd4075;
          lut[8081] <= 16'd4318;
          lut[8082] <= 16'd4560;
          lut[8083] <= 16'd4799;
          lut[8084] <= 16'd5036;
          lut[8085] <= 16'd5272;
          lut[8086] <= 16'd5504;
          lut[8087] <= 16'd5735;
          lut[8088] <= 16'd5963;
          lut[8089] <= 16'd6189;
          lut[8090] <= 16'd6413;
          lut[8091] <= 16'd6634;
          lut[8092] <= 16'd6852;
          lut[8093] <= 16'd7068;
          lut[8094] <= 16'd7281;
          lut[8095] <= 16'd7492;
          lut[8096] <= 16'd7700;
          lut[8097] <= 16'd7905;
          lut[8098] <= 16'd8108;
          lut[8099] <= 16'd8308;
          lut[8100] <= 16'd8506;
          lut[8101] <= 16'd8700;
          lut[8102] <= 16'd8892;
          lut[8103] <= 16'd9082;
          lut[8104] <= 16'd9268;
          lut[8105] <= 16'd9452;
          lut[8106] <= 16'd9634;
          lut[8107] <= 16'd9813;
          lut[8108] <= 16'd9989;
          lut[8109] <= 16'd10162;
          lut[8110] <= 16'd10333;
          lut[8111] <= 16'd10501;
          lut[8112] <= 16'd10667;
          lut[8113] <= 16'd10831;
          lut[8114] <= 16'd10991;
          lut[8115] <= 16'd11150;
          lut[8116] <= 16'd11306;
          lut[8117] <= 16'd11459;
          lut[8118] <= 16'd11610;
          lut[8119] <= 16'd11759;
          lut[8120] <= 16'd11905;
          lut[8121] <= 16'd12049;
          lut[8122] <= 16'd12191;
          lut[8123] <= 16'd12331;
          lut[8124] <= 16'd12468;
          lut[8125] <= 16'd12604;
          lut[8126] <= 16'd12737;
          lut[8127] <= 16'd12868;
          lut[8128] <= 16'd12997;
          lut[8129] <= 16'd13124;
          lut[8130] <= 16'd13249;
          lut[8131] <= 16'd13372;
          lut[8132] <= 16'd13493;
          lut[8133] <= 16'd13612;
          lut[8134] <= 16'd13729;
          lut[8135] <= 16'd13845;
          lut[8136] <= 16'd13959;
          lut[8137] <= 16'd14071;
          lut[8138] <= 16'd14181;
          lut[8139] <= 16'd14289;
          lut[8140] <= 16'd14396;
          lut[8141] <= 16'd14501;
          lut[8142] <= 16'd14604;
          lut[8143] <= 16'd14706;
          lut[8144] <= 16'd14807;
          lut[8145] <= 16'd14905;
          lut[8146] <= 16'd15003;
          lut[8147] <= 16'd15098;
          lut[8148] <= 16'd15193;
          lut[8149] <= 16'd15286;
          lut[8150] <= 16'd15377;
          lut[8151] <= 16'd15467;
          lut[8152] <= 16'd15556;
          lut[8153] <= 16'd15644;
          lut[8154] <= 16'd15730;
          lut[8155] <= 16'd15815;
          lut[8156] <= 16'd15898;
          lut[8157] <= 16'd15981;
          lut[8158] <= 16'd16062;
          lut[8159] <= 16'd16142;
          lut[8160] <= 16'd16221;
          lut[8161] <= 16'd16299;
          lut[8162] <= 16'd16375;
          lut[8163] <= 16'd16451;
          lut[8164] <= 16'd16525;
          lut[8165] <= 16'd16598;
          lut[8166] <= 16'd16671;
          lut[8167] <= 16'd16742;
          lut[8168] <= 16'd16812;
          lut[8169] <= 16'd16882;
          lut[8170] <= 16'd16950;
          lut[8171] <= 16'd17017;
          lut[8172] <= 16'd17084;
          lut[8173] <= 16'd17150;
          lut[8174] <= 16'd17214;
          lut[8175] <= 16'd17278;
          lut[8176] <= 16'd17341;
          lut[8177] <= 16'd17403;
          lut[8178] <= 16'd17464;
          lut[8179] <= 16'd17525;
          lut[8180] <= 16'd17584;
          lut[8181] <= 16'd17643;
          lut[8182] <= 16'd17701;
          lut[8183] <= 16'd17759;
          lut[8184] <= 16'd17815;
          lut[8185] <= 16'd17871;
          lut[8186] <= 16'd17926;
          lut[8187] <= 16'd17980;
          lut[8188] <= 16'd18034;
          lut[8189] <= 16'd18087;
          lut[8190] <= 16'd18140;
          lut[8191] <= 16'd18191;
          lut[8192] <= 0;
          lut[8193] <= 16'd256;
          lut[8194] <= 16'd512;
          lut[8195] <= 16'd767;
          lut[8196] <= 16'd1023;
          lut[8197] <= 16'd1277;
          lut[8198] <= 16'd1532;
          lut[8199] <= 16'd1785;
          lut[8200] <= 16'd2037;
          lut[8201] <= 16'd2289;
          lut[8202] <= 16'd2539;
          lut[8203] <= 16'd2789;
          lut[8204] <= 16'd3037;
          lut[8205] <= 16'd3283;
          lut[8206] <= 16'd3528;
          lut[8207] <= 16'd3772;
          lut[8208] <= 16'd4014;
          lut[8209] <= 16'd4254;
          lut[8210] <= 16'd4492;
          lut[8211] <= 16'd4728;
          lut[8212] <= 16'd4962;
          lut[8213] <= 16'd5195;
          lut[8214] <= 16'd5425;
          lut[8215] <= 16'd5653;
          lut[8216] <= 16'd5878;
          lut[8217] <= 16'd6101;
          lut[8218] <= 16'd6322;
          lut[8219] <= 16'd6541;
          lut[8220] <= 16'd6757;
          lut[8221] <= 16'd6971;
          lut[8222] <= 16'd7182;
          lut[8223] <= 16'd7390;
          lut[8224] <= 16'd7596;
          lut[8225] <= 16'd7800;
          lut[8226] <= 16'd8001;
          lut[8227] <= 16'd8199;
          lut[8228] <= 16'd8395;
          lut[8229] <= 16'd8588;
          lut[8230] <= 16'd8779;
          lut[8231] <= 16'd8967;
          lut[8232] <= 16'd9152;
          lut[8233] <= 16'd9335;
          lut[8234] <= 16'd9515;
          lut[8235] <= 16'd9693;
          lut[8236] <= 16'd9868;
          lut[8237] <= 16'd10040;
          lut[8238] <= 16'd10210;
          lut[8239] <= 16'd10378;
          lut[8240] <= 16'd10543;
          lut[8241] <= 16'd10706;
          lut[8242] <= 16'd10866;
          lut[8243] <= 16'd11024;
          lut[8244] <= 16'd11179;
          lut[8245] <= 16'd11332;
          lut[8246] <= 16'd11483;
          lut[8247] <= 16'd11631;
          lut[8248] <= 16'd11777;
          lut[8249] <= 16'd11921;
          lut[8250] <= 16'd12063;
          lut[8251] <= 16'd12202;
          lut[8252] <= 16'd12340;
          lut[8253] <= 16'd12475;
          lut[8254] <= 16'd12608;
          lut[8255] <= 16'd12739;
          lut[8256] <= 16'd12868;
          lut[8257] <= 16'd12995;
          lut[8258] <= 16'd13120;
          lut[8259] <= 16'd13243;
          lut[8260] <= 16'd13364;
          lut[8261] <= 16'd13484;
          lut[8262] <= 16'd13601;
          lut[8263] <= 16'd13717;
          lut[8264] <= 16'd13831;
          lut[8265] <= 16'd13943;
          lut[8266] <= 16'd14053;
          lut[8267] <= 16'd14162;
          lut[8268] <= 16'd14269;
          lut[8269] <= 16'd14374;
          lut[8270] <= 16'd14478;
          lut[8271] <= 16'd14580;
          lut[8272] <= 16'd14681;
          lut[8273] <= 16'd14780;
          lut[8274] <= 16'd14878;
          lut[8275] <= 16'd14974;
          lut[8276] <= 16'd15069;
          lut[8277] <= 16'd15162;
          lut[8278] <= 16'd15254;
          lut[8279] <= 16'd15345;
          lut[8280] <= 16'd15434;
          lut[8281] <= 16'd15522;
          lut[8282] <= 16'd15608;
          lut[8283] <= 16'd15694;
          lut[8284] <= 16'd15778;
          lut[8285] <= 16'd15861;
          lut[8286] <= 16'd15942;
          lut[8287] <= 16'd16023;
          lut[8288] <= 16'd16102;
          lut[8289] <= 16'd16180;
          lut[8290] <= 16'd16257;
          lut[8291] <= 16'd16333;
          lut[8292] <= 16'd16408;
          lut[8293] <= 16'd16482;
          lut[8294] <= 16'd16555;
          lut[8295] <= 16'd16627;
          lut[8296] <= 16'd16698;
          lut[8297] <= 16'd16767;
          lut[8298] <= 16'd16836;
          lut[8299] <= 16'd16904;
          lut[8300] <= 16'd16971;
          lut[8301] <= 16'd17037;
          lut[8302] <= 16'd17102;
          lut[8303] <= 16'd17167;
          lut[8304] <= 16'd17230;
          lut[8305] <= 16'd17293;
          lut[8306] <= 16'd17355;
          lut[8307] <= 16'd17416;
          lut[8308] <= 16'd17476;
          lut[8309] <= 16'd17535;
          lut[8310] <= 16'd17594;
          lut[8311] <= 16'd17651;
          lut[8312] <= 16'd17708;
          lut[8313] <= 16'd17765;
          lut[8314] <= 16'd17820;
          lut[8315] <= 16'd17875;
          lut[8316] <= 16'd17929;
          lut[8317] <= 16'd17983;
          lut[8318] <= 16'd18036;
          lut[8319] <= 16'd18088;
          lut[8320] <= 0;
          lut[8321] <= 16'd252;
          lut[8322] <= 16'd504;
          lut[8323] <= 16'd756;
          lut[8324] <= 16'd1007;
          lut[8325] <= 16'd1258;
          lut[8326] <= 16'd1508;
          lut[8327] <= 16'd1758;
          lut[8328] <= 16'd2006;
          lut[8329] <= 16'd2254;
          lut[8330] <= 16'd2501;
          lut[8331] <= 16'd2747;
          lut[8332] <= 16'd2991;
          lut[8333] <= 16'd3234;
          lut[8334] <= 16'd3476;
          lut[8335] <= 16'd3716;
          lut[8336] <= 16'd3954;
          lut[8337] <= 16'd4191;
          lut[8338] <= 16'd4426;
          lut[8339] <= 16'd4659;
          lut[8340] <= 16'd4891;
          lut[8341] <= 16'd5120;
          lut[8342] <= 16'd5347;
          lut[8343] <= 16'd5572;
          lut[8344] <= 16'd5795;
          lut[8345] <= 16'd6016;
          lut[8346] <= 16'd6234;
          lut[8347] <= 16'd6450;
          lut[8348] <= 16'd6664;
          lut[8349] <= 16'd6876;
          lut[8350] <= 16'd7085;
          lut[8351] <= 16'd7291;
          lut[8352] <= 16'd7495;
          lut[8353] <= 16'd7697;
          lut[8354] <= 16'd7896;
          lut[8355] <= 16'd8093;
          lut[8356] <= 16'd8287;
          lut[8357] <= 16'd8479;
          lut[8358] <= 16'd8668;
          lut[8359] <= 16'd8854;
          lut[8360] <= 16'd9038;
          lut[8361] <= 16'd9220;
          lut[8362] <= 16'd9399;
          lut[8363] <= 16'd9576;
          lut[8364] <= 16'd9750;
          lut[8365] <= 16'd9921;
          lut[8366] <= 16'd10090;
          lut[8367] <= 16'd10257;
          lut[8368] <= 16'd10421;
          lut[8369] <= 16'd10583;
          lut[8370] <= 16'd10743;
          lut[8371] <= 16'd10900;
          lut[8372] <= 16'd11055;
          lut[8373] <= 16'd11208;
          lut[8374] <= 16'd11358;
          lut[8375] <= 16'd11506;
          lut[8376] <= 16'd11652;
          lut[8377] <= 16'd11795;
          lut[8378] <= 16'd11937;
          lut[8379] <= 16'd12076;
          lut[8380] <= 16'd12213;
          lut[8381] <= 16'd12348;
          lut[8382] <= 16'd12481;
          lut[8383] <= 16'd12612;
          lut[8384] <= 16'd12741;
          lut[8385] <= 16'd12868;
          lut[8386] <= 16'd12993;
          lut[8387] <= 16'd13116;
          lut[8388] <= 16'd13237;
          lut[8389] <= 16'd13357;
          lut[8390] <= 16'd13475;
          lut[8391] <= 16'd13590;
          lut[8392] <= 16'd13704;
          lut[8393] <= 16'd13817;
          lut[8394] <= 16'd13927;
          lut[8395] <= 16'd14036;
          lut[8396] <= 16'd14144;
          lut[8397] <= 16'd14249;
          lut[8398] <= 16'd14353;
          lut[8399] <= 16'd14456;
          lut[8400] <= 16'd14557;
          lut[8401] <= 16'd14656;
          lut[8402] <= 16'd14754;
          lut[8403] <= 16'd14851;
          lut[8404] <= 16'd14946;
          lut[8405] <= 16'd15040;
          lut[8406] <= 16'd15132;
          lut[8407] <= 16'd15223;
          lut[8408] <= 16'd15313;
          lut[8409] <= 16'd15401;
          lut[8410] <= 16'd15488;
          lut[8411] <= 16'd15574;
          lut[8412] <= 16'd15658;
          lut[8413] <= 16'd15742;
          lut[8414] <= 16'd15824;
          lut[8415] <= 16'd15905;
          lut[8416] <= 16'd15985;
          lut[8417] <= 16'd16063;
          lut[8418] <= 16'd16141;
          lut[8419] <= 16'd16217;
          lut[8420] <= 16'd16293;
          lut[8421] <= 16'd16367;
          lut[8422] <= 16'd16440;
          lut[8423] <= 16'd16513;
          lut[8424] <= 16'd16584;
          lut[8425] <= 16'd16654;
          lut[8426] <= 16'd16724;
          lut[8427] <= 16'd16792;
          lut[8428] <= 16'd16859;
          lut[8429] <= 16'd16926;
          lut[8430] <= 16'd16992;
          lut[8431] <= 16'd17056;
          lut[8432] <= 16'd17120;
          lut[8433] <= 16'd17183;
          lut[8434] <= 16'd17246;
          lut[8435] <= 16'd17307;
          lut[8436] <= 16'd17368;
          lut[8437] <= 16'd17428;
          lut[8438] <= 16'd17487;
          lut[8439] <= 16'd17545;
          lut[8440] <= 16'd17603;
          lut[8441] <= 16'd17659;
          lut[8442] <= 16'd17715;
          lut[8443] <= 16'd17771;
          lut[8444] <= 16'd17825;
          lut[8445] <= 16'd17879;
          lut[8446] <= 16'd17933;
          lut[8447] <= 16'd17985;
          lut[8448] <= 0;
          lut[8449] <= 16'd248;
          lut[8450] <= 16'd496;
          lut[8451] <= 16'd744;
          lut[8452] <= 16'd992;
          lut[8453] <= 16'd1239;
          lut[8454] <= 16'd1485;
          lut[8455] <= 16'd1731;
          lut[8456] <= 16'd1976;
          lut[8457] <= 16'd2220;
          lut[8458] <= 16'd2464;
          lut[8459] <= 16'd2706;
          lut[8460] <= 16'd2947;
          lut[8461] <= 16'd3186;
          lut[8462] <= 16'd3425;
          lut[8463] <= 16'd3661;
          lut[8464] <= 16'd3897;
          lut[8465] <= 16'd4130;
          lut[8466] <= 16'd4362;
          lut[8467] <= 16'd4592;
          lut[8468] <= 16'd4821;
          lut[8469] <= 16'd5047;
          lut[8470] <= 16'd5272;
          lut[8471] <= 16'd5494;
          lut[8472] <= 16'd5714;
          lut[8473] <= 16'd5932;
          lut[8474] <= 16'd6148;
          lut[8475] <= 16'd6362;
          lut[8476] <= 16'd6574;
          lut[8477] <= 16'd6783;
          lut[8478] <= 16'd6990;
          lut[8479] <= 16'd7194;
          lut[8480] <= 16'd7397;
          lut[8481] <= 16'd7596;
          lut[8482] <= 16'd7794;
          lut[8483] <= 16'd7989;
          lut[8484] <= 16'd8181;
          lut[8485] <= 16'd8371;
          lut[8486] <= 16'd8559;
          lut[8487] <= 16'd8744;
          lut[8488] <= 16'd8927;
          lut[8489] <= 16'd9107;
          lut[8490] <= 16'd9285;
          lut[8491] <= 16'd9461;
          lut[8492] <= 16'd9634;
          lut[8493] <= 16'd9804;
          lut[8494] <= 16'd9973;
          lut[8495] <= 16'd10139;
          lut[8496] <= 16'd10302;
          lut[8497] <= 16'd10463;
          lut[8498] <= 16'd10622;
          lut[8499] <= 16'd10779;
          lut[8500] <= 16'd10933;
          lut[8501] <= 16'd11085;
          lut[8502] <= 16'd11235;
          lut[8503] <= 16'd11383;
          lut[8504] <= 16'd11528;
          lut[8505] <= 16'd11671;
          lut[8506] <= 16'd11812;
          lut[8507] <= 16'd11951;
          lut[8508] <= 16'd12088;
          lut[8509] <= 16'd12223;
          lut[8510] <= 16'd12356;
          lut[8511] <= 16'd12487;
          lut[8512] <= 16'd12616;
          lut[8513] <= 16'd12743;
          lut[8514] <= 16'd12868;
          lut[8515] <= 16'd12991;
          lut[8516] <= 16'd13112;
          lut[8517] <= 16'd13232;
          lut[8518] <= 16'd13350;
          lut[8519] <= 16'd13466;
          lut[8520] <= 16'd13580;
          lut[8521] <= 16'd13692;
          lut[8522] <= 16'd13803;
          lut[8523] <= 16'd13912;
          lut[8524] <= 16'd14020;
          lut[8525] <= 16'd14126;
          lut[8526] <= 16'd14230;
          lut[8527] <= 16'd14333;
          lut[8528] <= 16'd14434;
          lut[8529] <= 16'd14534;
          lut[8530] <= 16'd14632;
          lut[8531] <= 16'd14729;
          lut[8532] <= 16'd14825;
          lut[8533] <= 16'd14919;
          lut[8534] <= 16'd15011;
          lut[8535] <= 16'd15103;
          lut[8536] <= 16'd15193;
          lut[8537] <= 16'd15282;
          lut[8538] <= 16'd15369;
          lut[8539] <= 16'd15455;
          lut[8540] <= 16'd15540;
          lut[8541] <= 16'd15624;
          lut[8542] <= 16'd15706;
          lut[8543] <= 16'd15788;
          lut[8544] <= 16'd15868;
          lut[8545] <= 16'd15947;
          lut[8546] <= 16'd16025;
          lut[8547] <= 16'd16102;
          lut[8548] <= 16'd16178;
          lut[8549] <= 16'd16253;
          lut[8550] <= 16'd16327;
          lut[8551] <= 16'd16399;
          lut[8552] <= 16'd16471;
          lut[8553] <= 16'd16542;
          lut[8554] <= 16'd16612;
          lut[8555] <= 16'd16681;
          lut[8556] <= 16'd16748;
          lut[8557] <= 16'd16816;
          lut[8558] <= 16'd16882;
          lut[8559] <= 16'd16947;
          lut[8560] <= 16'd17011;
          lut[8561] <= 16'd17075;
          lut[8562] <= 16'd17138;
          lut[8563] <= 16'd17200;
          lut[8564] <= 16'd17261;
          lut[8565] <= 16'd17321;
          lut[8566] <= 16'd17381;
          lut[8567] <= 16'd17439;
          lut[8568] <= 16'd17497;
          lut[8569] <= 16'd17555;
          lut[8570] <= 16'd17611;
          lut[8571] <= 16'd17667;
          lut[8572] <= 16'd17722;
          lut[8573] <= 16'd17777;
          lut[8574] <= 16'd17830;
          lut[8575] <= 16'd17884;
          lut[8576] <= 0;
          lut[8577] <= 16'd245;
          lut[8578] <= 16'd489;
          lut[8579] <= 16'd733;
          lut[8580] <= 16'd977;
          lut[8581] <= 16'd1220;
          lut[8582] <= 16'd1463;
          lut[8583] <= 16'd1706;
          lut[8584] <= 16'd1947;
          lut[8585] <= 16'd2188;
          lut[8586] <= 16'd2427;
          lut[8587] <= 16'd2666;
          lut[8588] <= 16'd2904;
          lut[8589] <= 16'd3140;
          lut[8590] <= 16'd3375;
          lut[8591] <= 16'd3609;
          lut[8592] <= 16'd3841;
          lut[8593] <= 16'd4071;
          lut[8594] <= 16'd4300;
          lut[8595] <= 16'd4527;
          lut[8596] <= 16'd4753;
          lut[8597] <= 16'd4976;
          lut[8598] <= 16'd5198;
          lut[8599] <= 16'd5418;
          lut[8600] <= 16'd5636;
          lut[8601] <= 16'd5851;
          lut[8602] <= 16'd6065;
          lut[8603] <= 16'd6276;
          lut[8604] <= 16'd6486;
          lut[8605] <= 16'd6693;
          lut[8606] <= 16'd6898;
          lut[8607] <= 16'd7100;
          lut[8608] <= 16'd7300;
          lut[8609] <= 16'd7498;
          lut[8610] <= 16'd7694;
          lut[8611] <= 16'd7887;
          lut[8612] <= 16'd8078;
          lut[8613] <= 16'd8267;
          lut[8614] <= 16'd8453;
          lut[8615] <= 16'd8637;
          lut[8616] <= 16'd8818;
          lut[8617] <= 16'd8997;
          lut[8618] <= 16'd9174;
          lut[8619] <= 16'd9348;
          lut[8620] <= 16'd9520;
          lut[8621] <= 16'd9690;
          lut[8622] <= 16'd9857;
          lut[8623] <= 16'd10023;
          lut[8624] <= 16'd10185;
          lut[8625] <= 16'd10346;
          lut[8626] <= 16'd10504;
          lut[8627] <= 16'd10660;
          lut[8628] <= 16'd10814;
          lut[8629] <= 16'd10965;
          lut[8630] <= 16'd11114;
          lut[8631] <= 16'd11262;
          lut[8632] <= 16'd11407;
          lut[8633] <= 16'd11550;
          lut[8634] <= 16'd11690;
          lut[8635] <= 16'd11829;
          lut[8636] <= 16'd11966;
          lut[8637] <= 16'd12101;
          lut[8638] <= 16'd12233;
          lut[8639] <= 16'd12364;
          lut[8640] <= 16'd12493;
          lut[8641] <= 16'd12620;
          lut[8642] <= 16'd12745;
          lut[8643] <= 16'd12868;
          lut[8644] <= 16'd12989;
          lut[8645] <= 16'd13109;
          lut[8646] <= 16'd13227;
          lut[8647] <= 16'd13343;
          lut[8648] <= 16'd13457;
          lut[8649] <= 16'd13570;
          lut[8650] <= 16'd13681;
          lut[8651] <= 16'd13790;
          lut[8652] <= 16'd13898;
          lut[8653] <= 16'd14004;
          lut[8654] <= 16'd14109;
          lut[8655] <= 16'd14212;
          lut[8656] <= 16'd14313;
          lut[8657] <= 16'd14413;
          lut[8658] <= 16'd14512;
          lut[8659] <= 16'd14609;
          lut[8660] <= 16'd14705;
          lut[8661] <= 16'd14799;
          lut[8662] <= 16'd14892;
          lut[8663] <= 16'd14984;
          lut[8664] <= 16'd15074;
          lut[8665] <= 16'd15163;
          lut[8666] <= 16'd15251;
          lut[8667] <= 16'd15338;
          lut[8668] <= 16'd15423;
          lut[8669] <= 16'd15507;
          lut[8670] <= 16'd15590;
          lut[8671] <= 16'd15672;
          lut[8672] <= 16'd15753;
          lut[8673] <= 16'd15832;
          lut[8674] <= 16'd15911;
          lut[8675] <= 16'd15988;
          lut[8676] <= 16'd16064;
          lut[8677] <= 16'd16140;
          lut[8678] <= 16'd16214;
          lut[8679] <= 16'd16287;
          lut[8680] <= 16'd16359;
          lut[8681] <= 16'd16430;
          lut[8682] <= 16'd16501;
          lut[8683] <= 16'd16570;
          lut[8684] <= 16'd16638;
          lut[8685] <= 16'd16706;
          lut[8686] <= 16'd16773;
          lut[8687] <= 16'd16838;
          lut[8688] <= 16'd16903;
          lut[8689] <= 16'd16967;
          lut[8690] <= 16'd17030;
          lut[8691] <= 16'd17093;
          lut[8692] <= 16'd17154;
          lut[8693] <= 16'd17215;
          lut[8694] <= 16'd17275;
          lut[8695] <= 16'd17334;
          lut[8696] <= 16'd17393;
          lut[8697] <= 16'd17451;
          lut[8698] <= 16'd17508;
          lut[8699] <= 16'd17564;
          lut[8700] <= 16'd17620;
          lut[8701] <= 16'd17674;
          lut[8702] <= 16'd17729;
          lut[8703] <= 16'd17782;
          lut[8704] <= 0;
          lut[8705] <= 16'd241;
          lut[8706] <= 16'd482;
          lut[8707] <= 16'd722;
          lut[8708] <= 16'd963;
          lut[8709] <= 16'd1203;
          lut[8710] <= 16'd1442;
          lut[8711] <= 16'd1681;
          lut[8712] <= 16'd1919;
          lut[8713] <= 16'd2156;
          lut[8714] <= 16'd2392;
          lut[8715] <= 16'd2628;
          lut[8716] <= 16'd2862;
          lut[8717] <= 16'd3095;
          lut[8718] <= 16'd3327;
          lut[8719] <= 16'd3557;
          lut[8720] <= 16'd3786;
          lut[8721] <= 16'd4014;
          lut[8722] <= 16'd4240;
          lut[8723] <= 16'd4464;
          lut[8724] <= 16'd4687;
          lut[8725] <= 16'd4908;
          lut[8726] <= 16'd5127;
          lut[8727] <= 16'd5344;
          lut[8728] <= 16'd5559;
          lut[8729] <= 16'd5772;
          lut[8730] <= 16'd5983;
          lut[8731] <= 16'd6193;
          lut[8732] <= 16'd6400;
          lut[8733] <= 16'd6605;
          lut[8734] <= 16'd6807;
          lut[8735] <= 16'd7008;
          lut[8736] <= 16'd7206;
          lut[8737] <= 16'd7403;
          lut[8738] <= 16'd7596;
          lut[8739] <= 16'd7788;
          lut[8740] <= 16'd7977;
          lut[8741] <= 16'd8164;
          lut[8742] <= 16'd8349;
          lut[8743] <= 16'd8532;
          lut[8744] <= 16'd8712;
          lut[8745] <= 16'd8890;
          lut[8746] <= 16'd9065;
          lut[8747] <= 16'd9238;
          lut[8748] <= 16'd9409;
          lut[8749] <= 16'd9578;
          lut[8750] <= 16'd9745;
          lut[8751] <= 16'd9909;
          lut[8752] <= 16'd10071;
          lut[8753] <= 16'd10230;
          lut[8754] <= 16'd10388;
          lut[8755] <= 16'd10543;
          lut[8756] <= 16'd10696;
          lut[8757] <= 16'd10847;
          lut[8758] <= 16'd10996;
          lut[8759] <= 16'd11143;
          lut[8760] <= 16'd11287;
          lut[8761] <= 16'd11430;
          lut[8762] <= 16'd11570;
          lut[8763] <= 16'd11709;
          lut[8764] <= 16'd11845;
          lut[8765] <= 16'd11980;
          lut[8766] <= 16'd12112;
          lut[8767] <= 16'd12243;
          lut[8768] <= 16'd12372;
          lut[8769] <= 16'd12498;
          lut[8770] <= 16'd12623;
          lut[8771] <= 16'd12747;
          lut[8772] <= 16'd12868;
          lut[8773] <= 16'd12988;
          lut[8774] <= 16'd13105;
          lut[8775] <= 16'd13222;
          lut[8776] <= 16'd13336;
          lut[8777] <= 16'd13449;
          lut[8778] <= 16'd13560;
          lut[8779] <= 16'd13669;
          lut[8780] <= 16'd13777;
          lut[8781] <= 16'd13884;
          lut[8782] <= 16'd13988;
          lut[8783] <= 16'd14092;
          lut[8784] <= 16'd14193;
          lut[8785] <= 16'd14294;
          lut[8786] <= 16'd14393;
          lut[8787] <= 16'd14490;
          lut[8788] <= 16'd14586;
          lut[8789] <= 16'd14681;
          lut[8790] <= 16'd14774;
          lut[8791] <= 16'd14866;
          lut[8792] <= 16'd14957;
          lut[8793] <= 16'd15047;
          lut[8794] <= 16'd15135;
          lut[8795] <= 16'd15222;
          lut[8796] <= 16'd15307;
          lut[8797] <= 16'd15392;
          lut[8798] <= 16'd15475;
          lut[8799] <= 16'd15557;
          lut[8800] <= 16'd15639;
          lut[8801] <= 16'd15718;
          lut[8802] <= 16'd15797;
          lut[8803] <= 16'd15875;
          lut[8804] <= 16'd15952;
          lut[8805] <= 16'd16027;
          lut[8806] <= 16'd16102;
          lut[8807] <= 16'd16176;
          lut[8808] <= 16'd16248;
          lut[8809] <= 16'd16320;
          lut[8810] <= 16'd16391;
          lut[8811] <= 16'd16461;
          lut[8812] <= 16'd16529;
          lut[8813] <= 16'd16597;
          lut[8814] <= 16'd16664;
          lut[8815] <= 16'd16731;
          lut[8816] <= 16'd16796;
          lut[8817] <= 16'd16860;
          lut[8818] <= 16'd16924;
          lut[8819] <= 16'd16987;
          lut[8820] <= 16'd17049;
          lut[8821] <= 16'd17110;
          lut[8822] <= 16'd17171;
          lut[8823] <= 16'd17230;
          lut[8824] <= 16'd17289;
          lut[8825] <= 16'd17347;
          lut[8826] <= 16'd17405;
          lut[8827] <= 16'd17462;
          lut[8828] <= 16'd17518;
          lut[8829] <= 16'd17573;
          lut[8830] <= 16'd17628;
          lut[8831] <= 16'd17682;
          lut[8832] <= 0;
          lut[8833] <= 16'd237;
          lut[8834] <= 16'd475;
          lut[8835] <= 16'd712;
          lut[8836] <= 16'd949;
          lut[8837] <= 16'd1185;
          lut[8838] <= 16'd1421;
          lut[8839] <= 16'd1656;
          lut[8840] <= 16'd1891;
          lut[8841] <= 16'd2125;
          lut[8842] <= 16'd2358;
          lut[8843] <= 16'd2590;
          lut[8844] <= 16'd2821;
          lut[8845] <= 16'd3051;
          lut[8846] <= 16'd3280;
          lut[8847] <= 16'd3507;
          lut[8848] <= 16'd3733;
          lut[8849] <= 16'd3958;
          lut[8850] <= 16'd4181;
          lut[8851] <= 16'd4402;
          lut[8852] <= 16'd4622;
          lut[8853] <= 16'd4841;
          lut[8854] <= 16'd5057;
          lut[8855] <= 16'd5272;
          lut[8856] <= 16'd5484;
          lut[8857] <= 16'd5695;
          lut[8858] <= 16'd5904;
          lut[8859] <= 16'd6111;
          lut[8860] <= 16'd6316;
          lut[8861] <= 16'd6519;
          lut[8862] <= 16'd6720;
          lut[8863] <= 16'd6918;
          lut[8864] <= 16'd7115;
          lut[8865] <= 16'd7309;
          lut[8866] <= 16'd7501;
          lut[8867] <= 16'd7691;
          lut[8868] <= 16'd7879;
          lut[8869] <= 16'd8064;
          lut[8870] <= 16'd8248;
          lut[8871] <= 16'd8429;
          lut[8872] <= 16'd8608;
          lut[8873] <= 16'd8784;
          lut[8874] <= 16'd8959;
          lut[8875] <= 16'd9131;
          lut[8876] <= 16'd9301;
          lut[8877] <= 16'd9468;
          lut[8878] <= 16'd9634;
          lut[8879] <= 16'd9797;
          lut[8880] <= 16'd9958;
          lut[8881] <= 16'd10117;
          lut[8882] <= 16'd10274;
          lut[8883] <= 16'd10429;
          lut[8884] <= 16'd10581;
          lut[8885] <= 16'd10731;
          lut[8886] <= 16'd10880;
          lut[8887] <= 16'd11026;
          lut[8888] <= 16'd11170;
          lut[8889] <= 16'd11312;
          lut[8890] <= 16'd11452;
          lut[8891] <= 16'd11591;
          lut[8892] <= 16'd11727;
          lut[8893] <= 16'd11861;
          lut[8894] <= 16'd11993;
          lut[8895] <= 16'd12124;
          lut[8896] <= 16'd12252;
          lut[8897] <= 16'd12379;
          lut[8898] <= 16'd12504;
          lut[8899] <= 16'd12627;
          lut[8900] <= 16'd12748;
          lut[8901] <= 16'd12868;
          lut[8902] <= 16'd12986;
          lut[8903] <= 16'd13102;
          lut[8904] <= 16'd13217;
          lut[8905] <= 16'd13329;
          lut[8906] <= 16'd13441;
          lut[8907] <= 16'd13550;
          lut[8908] <= 16'd13658;
          lut[8909] <= 16'd13765;
          lut[8910] <= 16'd13870;
          lut[8911] <= 16'd13973;
          lut[8912] <= 16'd14075;
          lut[8913] <= 16'd14176;
          lut[8914] <= 16'd14275;
          lut[8915] <= 16'd14373;
          lut[8916] <= 16'd14469;
          lut[8917] <= 16'd14564;
          lut[8918] <= 16'd14658;
          lut[8919] <= 16'd14750;
          lut[8920] <= 16'd14841;
          lut[8921] <= 16'd14931;
          lut[8922] <= 16'd15019;
          lut[8923] <= 16'd15107;
          lut[8924] <= 16'd15193;
          lut[8925] <= 16'd15278;
          lut[8926] <= 16'd15361;
          lut[8927] <= 16'd15444;
          lut[8928] <= 16'd15525;
          lut[8929] <= 16'd15606;
          lut[8930] <= 16'd15685;
          lut[8931] <= 16'd15763;
          lut[8932] <= 16'd15840;
          lut[8933] <= 16'd15916;
          lut[8934] <= 16'd15991;
          lut[8935] <= 16'd16065;
          lut[8936] <= 16'd16139;
          lut[8937] <= 16'd16211;
          lut[8938] <= 16'd16282;
          lut[8939] <= 16'd16352;
          lut[8940] <= 16'd16421;
          lut[8941] <= 16'd16490;
          lut[8942] <= 16'd16557;
          lut[8943] <= 16'd16624;
          lut[8944] <= 16'd16689;
          lut[8945] <= 16'd16754;
          lut[8946] <= 16'd16818;
          lut[8947] <= 16'd16882;
          lut[8948] <= 16'd16944;
          lut[8949] <= 16'd17006;
          lut[8950] <= 16'd17067;
          lut[8951] <= 16'd17127;
          lut[8952] <= 16'd17186;
          lut[8953] <= 16'd17245;
          lut[8954] <= 16'd17303;
          lut[8955] <= 16'd17360;
          lut[8956] <= 16'd17416;
          lut[8957] <= 16'd17472;
          lut[8958] <= 16'd17527;
          lut[8959] <= 16'd17582;
          lut[8960] <= 0;
          lut[8961] <= 16'd234;
          lut[8962] <= 16'd468;
          lut[8963] <= 16'd702;
          lut[8964] <= 16'd935;
          lut[8965] <= 16'd1168;
          lut[8966] <= 16'd1401;
          lut[8967] <= 16'd1633;
          lut[8968] <= 16'd1864;
          lut[8969] <= 16'd2095;
          lut[8970] <= 16'd2325;
          lut[8971] <= 16'd2554;
          lut[8972] <= 16'd2782;
          lut[8973] <= 16'd3008;
          lut[8974] <= 16'd3234;
          lut[8975] <= 16'd3459;
          lut[8976] <= 16'd3682;
          lut[8977] <= 16'd3903;
          lut[8978] <= 16'd4124;
          lut[8979] <= 16'd4342;
          lut[8980] <= 16'd4560;
          lut[8981] <= 16'd4775;
          lut[8982] <= 16'd4989;
          lut[8983] <= 16'd5201;
          lut[8984] <= 16'd5412;
          lut[8985] <= 16'd5620;
          lut[8986] <= 16'd5827;
          lut[8987] <= 16'd6031;
          lut[8988] <= 16'd6234;
          lut[8989] <= 16'd6435;
          lut[8990] <= 16'd6634;
          lut[8991] <= 16'd6830;
          lut[8992] <= 16'd7025;
          lut[8993] <= 16'd7218;
          lut[8994] <= 16'd7408;
          lut[8995] <= 16'd7596;
          lut[8996] <= 16'd7783;
          lut[8997] <= 16'd7967;
          lut[8998] <= 16'd8148;
          lut[8999] <= 16'd8328;
          lut[9000] <= 16'd8506;
          lut[9001] <= 16'd8681;
          lut[9002] <= 16'd8854;
          lut[9003] <= 16'd9025;
          lut[9004] <= 16'd9194;
          lut[9005] <= 16'd9361;
          lut[9006] <= 16'd9525;
          lut[9007] <= 16'd9688;
          lut[9008] <= 16'd9848;
          lut[9009] <= 16'd10006;
          lut[9010] <= 16'd10162;
          lut[9011] <= 16'd10316;
          lut[9012] <= 16'd10468;
          lut[9013] <= 16'd10618;
          lut[9014] <= 16'd10766;
          lut[9015] <= 16'd10911;
          lut[9016] <= 16'd11055;
          lut[9017] <= 16'd11197;
          lut[9018] <= 16'd11336;
          lut[9019] <= 16'd11474;
          lut[9020] <= 16'd11610;
          lut[9021] <= 16'd11744;
          lut[9022] <= 16'd11876;
          lut[9023] <= 16'd12006;
          lut[9024] <= 16'd12135;
          lut[9025] <= 16'd12261;
          lut[9026] <= 16'd12386;
          lut[9027] <= 16'd12509;
          lut[9028] <= 16'd12631;
          lut[9029] <= 16'd12750;
          lut[9030] <= 16'd12868;
          lut[9031] <= 16'd12984;
          lut[9032] <= 16'd13099;
          lut[9033] <= 16'd13212;
          lut[9034] <= 16'd13323;
          lut[9035] <= 16'd13433;
          lut[9036] <= 16'd13541;
          lut[9037] <= 16'd13648;
          lut[9038] <= 16'd13753;
          lut[9039] <= 16'd13856;
          lut[9040] <= 16'd13959;
          lut[9041] <= 16'd14059;
          lut[9042] <= 16'd14159;
          lut[9043] <= 16'd14257;
          lut[9044] <= 16'd14353;
          lut[9045] <= 16'd14449;
          lut[9046] <= 16'd14543;
          lut[9047] <= 16'd14635;
          lut[9048] <= 16'd14726;
          lut[9049] <= 16'd14817;
          lut[9050] <= 16'd14905;
          lut[9051] <= 16'd14993;
          lut[9052] <= 16'd15079;
          lut[9053] <= 16'd15165;
          lut[9054] <= 16'd15249;
          lut[9055] <= 16'd15332;
          lut[9056] <= 16'd15413;
          lut[9057] <= 16'd15494;
          lut[9058] <= 16'd15574;
          lut[9059] <= 16'd15652;
          lut[9060] <= 16'd15730;
          lut[9061] <= 16'd15806;
          lut[9062] <= 16'd15882;
          lut[9063] <= 16'd15956;
          lut[9064] <= 16'd16030;
          lut[9065] <= 16'd16102;
          lut[9066] <= 16'd16174;
          lut[9067] <= 16'd16244;
          lut[9068] <= 16'd16314;
          lut[9069] <= 16'd16383;
          lut[9070] <= 16'd16451;
          lut[9071] <= 16'd16518;
          lut[9072] <= 16'd16584;
          lut[9073] <= 16'd16649;
          lut[9074] <= 16'd16714;
          lut[9075] <= 16'd16777;
          lut[9076] <= 16'd16840;
          lut[9077] <= 16'd16902;
          lut[9078] <= 16'd16964;
          lut[9079] <= 16'd17024;
          lut[9080] <= 16'd17084;
          lut[9081] <= 16'd17143;
          lut[9082] <= 16'd17201;
          lut[9083] <= 16'd17259;
          lut[9084] <= 16'd17316;
          lut[9085] <= 16'd17372;
          lut[9086] <= 16'd17428;
          lut[9087] <= 16'd17482;
          lut[9088] <= 0;
          lut[9089] <= 16'd231;
          lut[9090] <= 16'd461;
          lut[9091] <= 16'd692;
          lut[9092] <= 16'd922;
          lut[9093] <= 16'd1152;
          lut[9094] <= 16'd1381;
          lut[9095] <= 16'd1610;
          lut[9096] <= 16'd1838;
          lut[9097] <= 16'd2066;
          lut[9098] <= 16'd2293;
          lut[9099] <= 16'd2518;
          lut[9100] <= 16'd2743;
          lut[9101] <= 16'd2967;
          lut[9102] <= 16'd3190;
          lut[9103] <= 16'd3411;
          lut[9104] <= 16'd3632;
          lut[9105] <= 16'd3850;
          lut[9106] <= 16'd4068;
          lut[9107] <= 16'd4284;
          lut[9108] <= 16'd4499;
          lut[9109] <= 16'd4712;
          lut[9110] <= 16'd4923;
          lut[9111] <= 16'd5133;
          lut[9112] <= 16'd5341;
          lut[9113] <= 16'd5547;
          lut[9114] <= 16'd5751;
          lut[9115] <= 16'd5954;
          lut[9116] <= 16'd6154;
          lut[9117] <= 16'd6353;
          lut[9118] <= 16'd6550;
          lut[9119] <= 16'd6745;
          lut[9120] <= 16'd6938;
          lut[9121] <= 16'd7128;
          lut[9122] <= 16'd7317;
          lut[9123] <= 16'd7504;
          lut[9124] <= 16'd7688;
          lut[9125] <= 16'd7871;
          lut[9126] <= 16'd8051;
          lut[9127] <= 16'd8230;
          lut[9128] <= 16'd8406;
          lut[9129] <= 16'd8580;
          lut[9130] <= 16'd8752;
          lut[9131] <= 16'd8922;
          lut[9132] <= 16'd9090;
          lut[9133] <= 16'd9255;
          lut[9134] <= 16'd9419;
          lut[9135] <= 16'd9580;
          lut[9136] <= 16'd9740;
          lut[9137] <= 16'd9897;
          lut[9138] <= 16'd10053;
          lut[9139] <= 16'd10206;
          lut[9140] <= 16'd10357;
          lut[9141] <= 16'd10506;
          lut[9142] <= 16'd10653;
          lut[9143] <= 16'd10799;
          lut[9144] <= 16'd10942;
          lut[9145] <= 16'd11083;
          lut[9146] <= 16'd11222;
          lut[9147] <= 16'd11360;
          lut[9148] <= 16'd11495;
          lut[9149] <= 16'd11629;
          lut[9150] <= 16'd11761;
          lut[9151] <= 16'd11891;
          lut[9152] <= 16'd12019;
          lut[9153] <= 16'd12146;
          lut[9154] <= 16'd12270;
          lut[9155] <= 16'd12393;
          lut[9156] <= 16'd12514;
          lut[9157] <= 16'd12634;
          lut[9158] <= 16'd12752;
          lut[9159] <= 16'd12868;
          lut[9160] <= 16'd12983;
          lut[9161] <= 16'd13096;
          lut[9162] <= 16'd13207;
          lut[9163] <= 16'd13317;
          lut[9164] <= 16'd13425;
          lut[9165] <= 16'd13532;
          lut[9166] <= 16'd13637;
          lut[9167] <= 16'd13741;
          lut[9168] <= 16'd13843;
          lut[9169] <= 16'd13944;
          lut[9170] <= 16'd14044;
          lut[9171] <= 16'd14142;
          lut[9172] <= 16'd14239;
          lut[9173] <= 16'd14334;
          lut[9174] <= 16'd14429;
          lut[9175] <= 16'd14521;
          lut[9176] <= 16'd14613;
          lut[9177] <= 16'd14703;
          lut[9178] <= 16'd14793;
          lut[9179] <= 16'd14880;
          lut[9180] <= 16'd14967;
          lut[9181] <= 16'd15053;
          lut[9182] <= 16'd15137;
          lut[9183] <= 16'd15220;
          lut[9184] <= 16'd15303;
          lut[9185] <= 16'd15384;
          lut[9186] <= 16'd15464;
          lut[9187] <= 16'd15542;
          lut[9188] <= 16'd15620;
          lut[9189] <= 16'd15697;
          lut[9190] <= 16'd15773;
          lut[9191] <= 16'd15848;
          lut[9192] <= 16'd15922;
          lut[9193] <= 16'd15995;
          lut[9194] <= 16'd16066;
          lut[9195] <= 16'd16137;
          lut[9196] <= 16'd16208;
          lut[9197] <= 16'd16277;
          lut[9198] <= 16'd16345;
          lut[9199] <= 16'd16412;
          lut[9200] <= 16'd16479;
          lut[9201] <= 16'd16545;
          lut[9202] <= 16'd16610;
          lut[9203] <= 16'd16674;
          lut[9204] <= 16'd16737;
          lut[9205] <= 16'd16800;
          lut[9206] <= 16'd16861;
          lut[9207] <= 16'd16922;
          lut[9208] <= 16'd16982;
          lut[9209] <= 16'd17042;
          lut[9210] <= 16'd17101;
          lut[9211] <= 16'd17159;
          lut[9212] <= 16'd17216;
          lut[9213] <= 16'd17273;
          lut[9214] <= 16'd17329;
          lut[9215] <= 16'd17384;
          lut[9216] <= 0;
          lut[9217] <= 16'd228;
          lut[9218] <= 16'd455;
          lut[9219] <= 16'd682;
          lut[9220] <= 16'd909;
          lut[9221] <= 16'd1136;
          lut[9222] <= 16'd1362;
          lut[9223] <= 16'd1588;
          lut[9224] <= 16'd1813;
          lut[9225] <= 16'd2037;
          lut[9226] <= 16'd2261;
          lut[9227] <= 16'd2484;
          lut[9228] <= 16'd2706;
          lut[9229] <= 16'd2927;
          lut[9230] <= 16'd3147;
          lut[9231] <= 16'd3365;
          lut[9232] <= 16'd3583;
          lut[9233] <= 16'd3799;
          lut[9234] <= 16'd4014;
          lut[9235] <= 16'd4227;
          lut[9236] <= 16'd4439;
          lut[9237] <= 16'd4650;
          lut[9238] <= 16'd4859;
          lut[9239] <= 16'd5066;
          lut[9240] <= 16'd5272;
          lut[9241] <= 16'd5476;
          lut[9242] <= 16'd5678;
          lut[9243] <= 16'd5878;
          lut[9244] <= 16'd6077;
          lut[9245] <= 16'd6273;
          lut[9246] <= 16'd6468;
          lut[9247] <= 16'd6661;
          lut[9248] <= 16'd6852;
          lut[9249] <= 16'd7041;
          lut[9250] <= 16'd7228;
          lut[9251] <= 16'd7413;
          lut[9252] <= 16'd7596;
          lut[9253] <= 16'd7777;
          lut[9254] <= 16'd7956;
          lut[9255] <= 16'd8133;
          lut[9256] <= 16'd8308;
          lut[9257] <= 16'd8481;
          lut[9258] <= 16'd8652;
          lut[9259] <= 16'd8821;
          lut[9260] <= 16'd8987;
          lut[9261] <= 16'd9152;
          lut[9262] <= 16'd9315;
          lut[9263] <= 16'd9475;
          lut[9264] <= 16'd9634;
          lut[9265] <= 16'd9790;
          lut[9266] <= 16'd9945;
          lut[9267] <= 16'd10097;
          lut[9268] <= 16'd10248;
          lut[9269] <= 16'd10397;
          lut[9270] <= 16'd10543;
          lut[9271] <= 16'd10688;
          lut[9272] <= 16'd10831;
          lut[9273] <= 16'd10971;
          lut[9274] <= 16'd11110;
          lut[9275] <= 16'd11247;
          lut[9276] <= 16'd11383;
          lut[9277] <= 16'd11516;
          lut[9278] <= 16'd11648;
          lut[9279] <= 16'd11777;
          lut[9280] <= 16'd11905;
          lut[9281] <= 16'd12032;
          lut[9282] <= 16'd12156;
          lut[9283] <= 16'd12279;
          lut[9284] <= 16'd12400;
          lut[9285] <= 16'd12519;
          lut[9286] <= 16'd12637;
          lut[9287] <= 16'd12753;
          lut[9288] <= 16'd12868;
          lut[9289] <= 16'd12981;
          lut[9290] <= 16'd13092;
          lut[9291] <= 16'd13202;
          lut[9292] <= 16'd13311;
          lut[9293] <= 16'd13418;
          lut[9294] <= 16'd13523;
          lut[9295] <= 16'd13627;
          lut[9296] <= 16'd13729;
          lut[9297] <= 16'd13831;
          lut[9298] <= 16'd13930;
          lut[9299] <= 16'd14029;
          lut[9300] <= 16'd14126;
          lut[9301] <= 16'd14222;
          lut[9302] <= 16'd14316;
          lut[9303] <= 16'd14409;
          lut[9304] <= 16'd14501;
          lut[9305] <= 16'd14592;
          lut[9306] <= 16'd14681;
          lut[9307] <= 16'd14769;
          lut[9308] <= 16'd14856;
          lut[9309] <= 16'd14942;
          lut[9310] <= 16'd15027;
          lut[9311] <= 16'd15110;
          lut[9312] <= 16'd15193;
          lut[9313] <= 16'd15274;
          lut[9314] <= 16'd15354;
          lut[9315] <= 16'd15434;
          lut[9316] <= 16'd15512;
          lut[9317] <= 16'd15589;
          lut[9318] <= 16'd15665;
          lut[9319] <= 16'd15740;
          lut[9320] <= 16'd15815;
          lut[9321] <= 16'd15888;
          lut[9322] <= 16'd15960;
          lut[9323] <= 16'd16032;
          lut[9324] <= 16'd16102;
          lut[9325] <= 16'd16172;
          lut[9326] <= 16'd16240;
          lut[9327] <= 16'd16308;
          lut[9328] <= 16'd16375;
          lut[9329] <= 16'd16441;
          lut[9330] <= 16'd16507;
          lut[9331] <= 16'd16571;
          lut[9332] <= 16'd16635;
          lut[9333] <= 16'd16698;
          lut[9334] <= 16'd16760;
          lut[9335] <= 16'd16821;
          lut[9336] <= 16'd16882;
          lut[9337] <= 16'd16942;
          lut[9338] <= 16'd17001;
          lut[9339] <= 16'd17059;
          lut[9340] <= 16'd17117;
          lut[9341] <= 16'd17174;
          lut[9342] <= 16'd17230;
          lut[9343] <= 16'd17286;
          lut[9344] <= 0;
          lut[9345] <= 16'd224;
          lut[9346] <= 16'd449;
          lut[9347] <= 16'd673;
          lut[9348] <= 16'd897;
          lut[9349] <= 16'd1120;
          lut[9350] <= 16'd1344;
          lut[9351] <= 16'd1566;
          lut[9352] <= 16'd1788;
          lut[9353] <= 16'd2010;
          lut[9354] <= 16'd2231;
          lut[9355] <= 16'd2450;
          lut[9356] <= 16'd2669;
          lut[9357] <= 16'd2887;
          lut[9358] <= 16'd3104;
          lut[9359] <= 16'd3320;
          lut[9360] <= 16'd3535;
          lut[9361] <= 16'd3749;
          lut[9362] <= 16'd3961;
          lut[9363] <= 16'd4172;
          lut[9364] <= 16'd4381;
          lut[9365] <= 16'd4589;
          lut[9366] <= 16'd4796;
          lut[9367] <= 16'd5001;
          lut[9368] <= 16'd5204;
          lut[9369] <= 16'd5406;
          lut[9370] <= 16'd5606;
          lut[9371] <= 16'd5804;
          lut[9372] <= 16'd6001;
          lut[9373] <= 16'd6195;
          lut[9374] <= 16'd6388;
          lut[9375] <= 16'd6579;
          lut[9376] <= 16'd6769;
          lut[9377] <= 16'd6956;
          lut[9378] <= 16'd7141;
          lut[9379] <= 16'd7325;
          lut[9380] <= 16'd7506;
          lut[9381] <= 16'd7686;
          lut[9382] <= 16'd7864;
          lut[9383] <= 16'd8039;
          lut[9384] <= 16'd8213;
          lut[9385] <= 16'd8384;
          lut[9386] <= 16'd8554;
          lut[9387] <= 16'd8722;
          lut[9388] <= 16'd8887;
          lut[9389] <= 16'd9051;
          lut[9390] <= 16'd9212;
          lut[9391] <= 16'd9372;
          lut[9392] <= 16'd9530;
          lut[9393] <= 16'd9686;
          lut[9394] <= 16'd9839;
          lut[9395] <= 16'd9991;
          lut[9396] <= 16'd10141;
          lut[9397] <= 16'd10289;
          lut[9398] <= 16'd10435;
          lut[9399] <= 16'd10579;
          lut[9400] <= 16'd10721;
          lut[9401] <= 16'd10862;
          lut[9402] <= 16'd11000;
          lut[9403] <= 16'd11137;
          lut[9404] <= 16'd11272;
          lut[9405] <= 16'd11405;
          lut[9406] <= 16'd11536;
          lut[9407] <= 16'd11665;
          lut[9408] <= 16'd11793;
          lut[9409] <= 16'd11919;
          lut[9410] <= 16'd12044;
          lut[9411] <= 16'd12166;
          lut[9412] <= 16'd12287;
          lut[9413] <= 16'd12407;
          lut[9414] <= 16'd12524;
          lut[9415] <= 16'd12640;
          lut[9416] <= 16'd12755;
          lut[9417] <= 16'd12868;
          lut[9418] <= 16'd12979;
          lut[9419] <= 16'd13089;
          lut[9420] <= 16'd13198;
          lut[9421] <= 16'd13305;
          lut[9422] <= 16'd13410;
          lut[9423] <= 16'd13514;
          lut[9424] <= 16'd13617;
          lut[9425] <= 16'd13718;
          lut[9426] <= 16'd13818;
          lut[9427] <= 16'd13917;
          lut[9428] <= 16'd14014;
          lut[9429] <= 16'd14110;
          lut[9430] <= 16'd14205;
          lut[9431] <= 16'd14298;
          lut[9432] <= 16'd14390;
          lut[9433] <= 16'd14481;
          lut[9434] <= 16'd14571;
          lut[9435] <= 16'd14659;
          lut[9436] <= 16'd14746;
          lut[9437] <= 16'd14832;
          lut[9438] <= 16'd14917;
          lut[9439] <= 16'd15001;
          lut[9440] <= 16'd15084;
          lut[9441] <= 16'd15166;
          lut[9442] <= 16'd15246;
          lut[9443] <= 16'd15326;
          lut[9444] <= 16'd15405;
          lut[9445] <= 16'd15482;
          lut[9446] <= 16'd15559;
          lut[9447] <= 16'd15634;
          lut[9448] <= 16'd15709;
          lut[9449] <= 16'd15782;
          lut[9450] <= 16'd15855;
          lut[9451] <= 16'd15927;
          lut[9452] <= 16'd15998;
          lut[9453] <= 16'd16067;
          lut[9454] <= 16'd16137;
          lut[9455] <= 16'd16205;
          lut[9456] <= 16'd16272;
          lut[9457] <= 16'd16339;
          lut[9458] <= 16'd16404;
          lut[9459] <= 16'd16469;
          lut[9460] <= 16'd16533;
          lut[9461] <= 16'd16596;
          lut[9462] <= 16'd16659;
          lut[9463] <= 16'd16721;
          lut[9464] <= 16'd16782;
          lut[9465] <= 16'd16842;
          lut[9466] <= 16'd16901;
          lut[9467] <= 16'd16960;
          lut[9468] <= 16'd17018;
          lut[9469] <= 16'd17076;
          lut[9470] <= 16'd17133;
          lut[9471] <= 16'd17189;
          lut[9472] <= 0;
          lut[9473] <= 16'd221;
          lut[9474] <= 16'd443;
          lut[9475] <= 16'd664;
          lut[9476] <= 16'd885;
          lut[9477] <= 16'd1105;
          lut[9478] <= 16'd1326;
          lut[9479] <= 16'd1545;
          lut[9480] <= 16'd1764;
          lut[9481] <= 16'd1983;
          lut[9482] <= 16'd2201;
          lut[9483] <= 16'd2418;
          lut[9484] <= 16'd2634;
          lut[9485] <= 16'd2849;
          lut[9486] <= 16'd3063;
          lut[9487] <= 16'd3277;
          lut[9488] <= 16'd3489;
          lut[9489] <= 16'd3700;
          lut[9490] <= 16'd3909;
          lut[9491] <= 16'd4118;
          lut[9492] <= 16'd4325;
          lut[9493] <= 16'd4530;
          lut[9494] <= 16'd4735;
          lut[9495] <= 16'd4937;
          lut[9496] <= 16'd5138;
          lut[9497] <= 16'd5338;
          lut[9498] <= 16'd5536;
          lut[9499] <= 16'd5732;
          lut[9500] <= 16'd5927;
          lut[9501] <= 16'd6119;
          lut[9502] <= 16'd6310;
          lut[9503] <= 16'd6500;
          lut[9504] <= 16'd6687;
          lut[9505] <= 16'd6873;
          lut[9506] <= 16'd7056;
          lut[9507] <= 16'd7238;
          lut[9508] <= 16'd7418;
          lut[9509] <= 16'd7596;
          lut[9510] <= 16'd7773;
          lut[9511] <= 16'd7947;
          lut[9512] <= 16'd8119;
          lut[9513] <= 16'd8289;
          lut[9514] <= 16'd8458;
          lut[9515] <= 16'd8624;
          lut[9516] <= 16'd8789;
          lut[9517] <= 16'd8952;
          lut[9518] <= 16'd9112;
          lut[9519] <= 16'd9271;
          lut[9520] <= 16'd9428;
          lut[9521] <= 16'd9583;
          lut[9522] <= 16'd9736;
          lut[9523] <= 16'd9887;
          lut[9524] <= 16'd10036;
          lut[9525] <= 16'd10183;
          lut[9526] <= 16'd10328;
          lut[9527] <= 16'd10472;
          lut[9528] <= 16'd10614;
          lut[9529] <= 16'd10754;
          lut[9530] <= 16'd10892;
          lut[9531] <= 16'd11028;
          lut[9532] <= 16'd11162;
          lut[9533] <= 16'd11295;
          lut[9534] <= 16'd11426;
          lut[9535] <= 16'd11555;
          lut[9536] <= 16'd11683;
          lut[9537] <= 16'd11809;
          lut[9538] <= 16'd11933;
          lut[9539] <= 16'd12055;
          lut[9540] <= 16'd12176;
          lut[9541] <= 16'd12295;
          lut[9542] <= 16'd12413;
          lut[9543] <= 16'd12529;
          lut[9544] <= 16'd12644;
          lut[9545] <= 16'd12757;
          lut[9546] <= 16'd12868;
          lut[9547] <= 16'd12978;
          lut[9548] <= 16'd13086;
          lut[9549] <= 16'd13193;
          lut[9550] <= 16'd13299;
          lut[9551] <= 16'd13403;
          lut[9552] <= 16'd13506;
          lut[9553] <= 16'd13607;
          lut[9554] <= 16'd13707;
          lut[9555] <= 16'd13806;
          lut[9556] <= 16'd13904;
          lut[9557] <= 16'd14000;
          lut[9558] <= 16'd14094;
          lut[9559] <= 16'd14188;
          lut[9560] <= 16'd14280;
          lut[9561] <= 16'd14371;
          lut[9562] <= 16'd14461;
          lut[9563] <= 16'd14550;
          lut[9564] <= 16'd14638;
          lut[9565] <= 16'd14724;
          lut[9566] <= 16'd14809;
          lut[9567] <= 16'd14893;
          lut[9568] <= 16'd14977;
          lut[9569] <= 16'd15059;
          lut[9570] <= 16'd15139;
          lut[9571] <= 16'd15219;
          lut[9572] <= 16'd15298;
          lut[9573] <= 16'd15376;
          lut[9574] <= 16'd15453;
          lut[9575] <= 16'd15529;
          lut[9576] <= 16'd15604;
          lut[9577] <= 16'd15678;
          lut[9578] <= 16'd15751;
          lut[9579] <= 16'd15823;
          lut[9580] <= 16'd15894;
          lut[9581] <= 16'd15964;
          lut[9582] <= 16'd16034;
          lut[9583] <= 16'd16102;
          lut[9584] <= 16'd16170;
          lut[9585] <= 16'd16237;
          lut[9586] <= 16'd16303;
          lut[9587] <= 16'd16368;
          lut[9588] <= 16'd16432;
          lut[9589] <= 16'd16496;
          lut[9590] <= 16'd16559;
          lut[9591] <= 16'd16621;
          lut[9592] <= 16'd16682;
          lut[9593] <= 16'd16743;
          lut[9594] <= 16'd16803;
          lut[9595] <= 16'd16862;
          lut[9596] <= 16'd16921;
          lut[9597] <= 16'd16978;
          lut[9598] <= 16'd17036;
          lut[9599] <= 16'd17092;
          lut[9600] <= 0;
          lut[9601] <= 16'd218;
          lut[9602] <= 16'd437;
          lut[9603] <= 16'd655;
          lut[9604] <= 16'd873;
          lut[9605] <= 16'd1091;
          lut[9606] <= 16'd1308;
          lut[9607] <= 16'd1525;
          lut[9608] <= 16'd1741;
          lut[9609] <= 16'd1957;
          lut[9610] <= 16'd2172;
          lut[9611] <= 16'd2386;
          lut[9612] <= 16'd2599;
          lut[9613] <= 16'd2812;
          lut[9614] <= 16'd3024;
          lut[9615] <= 16'd3234;
          lut[9616] <= 16'd3444;
          lut[9617] <= 16'd3652;
          lut[9618] <= 16'd3859;
          lut[9619] <= 16'd4065;
          lut[9620] <= 16'd4270;
          lut[9621] <= 16'd4473;
          lut[9622] <= 16'd4675;
          lut[9623] <= 16'd4875;
          lut[9624] <= 16'd5074;
          lut[9625] <= 16'd5272;
          lut[9626] <= 16'd5467;
          lut[9627] <= 16'd5662;
          lut[9628] <= 16'd5854;
          lut[9629] <= 16'd6045;
          lut[9630] <= 16'd6234;
          lut[9631] <= 16'd6422;
          lut[9632] <= 16'd6607;
          lut[9633] <= 16'd6791;
          lut[9634] <= 16'd6973;
          lut[9635] <= 16'd7154;
          lut[9636] <= 16'd7332;
          lut[9637] <= 16'd7509;
          lut[9638] <= 16'd7684;
          lut[9639] <= 16'd7856;
          lut[9640] <= 16'd8027;
          lut[9641] <= 16'd8197;
          lut[9642] <= 16'd8364;
          lut[9643] <= 16'd8529;
          lut[9644] <= 16'd8693;
          lut[9645] <= 16'd8854;
          lut[9646] <= 16'd9014;
          lut[9647] <= 16'd9172;
          lut[9648] <= 16'd9328;
          lut[9649] <= 16'd9482;
          lut[9650] <= 16'd9634;
          lut[9651] <= 16'd9784;
          lut[9652] <= 16'd9933;
          lut[9653] <= 16'd10079;
          lut[9654] <= 16'd10224;
          lut[9655] <= 16'd10367;
          lut[9656] <= 16'd10508;
          lut[9657] <= 16'd10647;
          lut[9658] <= 16'd10785;
          lut[9659] <= 16'd10921;
          lut[9660] <= 16'd11055;
          lut[9661] <= 16'd11187;
          lut[9662] <= 16'd11318;
          lut[9663] <= 16'd11447;
          lut[9664] <= 16'd11574;
          lut[9665] <= 16'd11700;
          lut[9666] <= 16'd11824;
          lut[9667] <= 16'd11946;
          lut[9668] <= 16'd12067;
          lut[9669] <= 16'd12186;
          lut[9670] <= 16'd12303;
          lut[9671] <= 16'd12419;
          lut[9672] <= 16'd12534;
          lut[9673] <= 16'd12647;
          lut[9674] <= 16'd12758;
          lut[9675] <= 16'd12868;
          lut[9676] <= 16'd12976;
          lut[9677] <= 16'd13084;
          lut[9678] <= 16'd13189;
          lut[9679] <= 16'd13293;
          lut[9680] <= 16'd13396;
          lut[9681] <= 16'd13498;
          lut[9682] <= 16'd13598;
          lut[9683] <= 16'd13697;
          lut[9684] <= 16'd13794;
          lut[9685] <= 16'd13891;
          lut[9686] <= 16'd13986;
          lut[9687] <= 16'd14079;
          lut[9688] <= 16'd14172;
          lut[9689] <= 16'd14263;
          lut[9690] <= 16'd14353;
          lut[9691] <= 16'd14442;
          lut[9692] <= 16'd14530;
          lut[9693] <= 16'd14617;
          lut[9694] <= 16'd14702;
          lut[9695] <= 16'd14787;
          lut[9696] <= 16'd14870;
          lut[9697] <= 16'd14952;
          lut[9698] <= 16'd15033;
          lut[9699] <= 16'd15114;
          lut[9700] <= 16'd15193;
          lut[9701] <= 16'd15271;
          lut[9702] <= 16'd15348;
          lut[9703] <= 16'd15424;
          lut[9704] <= 16'd15499;
          lut[9705] <= 16'd15574;
          lut[9706] <= 16'd15647;
          lut[9707] <= 16'd15720;
          lut[9708] <= 16'd15791;
          lut[9709] <= 16'd15862;
          lut[9710] <= 16'd15931;
          lut[9711] <= 16'd16000;
          lut[9712] <= 16'd16068;
          lut[9713] <= 16'd16136;
          lut[9714] <= 16'd16202;
          lut[9715] <= 16'd16268;
          lut[9716] <= 16'd16332;
          lut[9717] <= 16'd16396;
          lut[9718] <= 16'd16460;
          lut[9719] <= 16'd16522;
          lut[9720] <= 16'd16584;
          lut[9721] <= 16'd16645;
          lut[9722] <= 16'd16705;
          lut[9723] <= 16'd16765;
          lut[9724] <= 16'd16824;
          lut[9725] <= 16'd16882;
          lut[9726] <= 16'd16939;
          lut[9727] <= 16'd16996;
          lut[9728] <= 0;
          lut[9729] <= 16'd216;
          lut[9730] <= 16'd431;
          lut[9731] <= 16'd646;
          lut[9732] <= 16'd862;
          lut[9733] <= 16'd1076;
          lut[9734] <= 16'd1291;
          lut[9735] <= 16'd1505;
          lut[9736] <= 16'd1718;
          lut[9737] <= 16'd1931;
          lut[9738] <= 16'd2143;
          lut[9739] <= 16'd2355;
          lut[9740] <= 16'd2566;
          lut[9741] <= 16'd2776;
          lut[9742] <= 16'd2985;
          lut[9743] <= 16'd3193;
          lut[9744] <= 16'd3400;
          lut[9745] <= 16'd3605;
          lut[9746] <= 16'd3810;
          lut[9747] <= 16'd4014;
          lut[9748] <= 16'd4216;
          lut[9749] <= 16'd4417;
          lut[9750] <= 16'd4617;
          lut[9751] <= 16'd4815;
          lut[9752] <= 16'd5012;
          lut[9753] <= 16'd5207;
          lut[9754] <= 16'd5401;
          lut[9755] <= 16'd5593;
          lut[9756] <= 16'd5783;
          lut[9757] <= 16'd5972;
          lut[9758] <= 16'd6160;
          lut[9759] <= 16'd6345;
          lut[9760] <= 16'd6529;
          lut[9761] <= 16'd6712;
          lut[9762] <= 16'd6892;
          lut[9763] <= 16'd7071;
          lut[9764] <= 16'd7248;
          lut[9765] <= 16'd7423;
          lut[9766] <= 16'd7596;
          lut[9767] <= 16'd7768;
          lut[9768] <= 16'd7938;
          lut[9769] <= 16'd8106;
          lut[9770] <= 16'd8272;
          lut[9771] <= 16'd8436;
          lut[9772] <= 16'd8598;
          lut[9773] <= 16'd8759;
          lut[9774] <= 16'd8917;
          lut[9775] <= 16'd9074;
          lut[9776] <= 16'd9229;
          lut[9777] <= 16'd9383;
          lut[9778] <= 16'd9534;
          lut[9779] <= 16'd9683;
          lut[9780] <= 16'd9831;
          lut[9781] <= 16'd9977;
          lut[9782] <= 16'd10121;
          lut[9783] <= 16'd10264;
          lut[9784] <= 16'd10404;
          lut[9785] <= 16'd10543;
          lut[9786] <= 16'd10680;
          lut[9787] <= 16'd10816;
          lut[9788] <= 16'd10949;
          lut[9789] <= 16'd11081;
          lut[9790] <= 16'd11211;
          lut[9791] <= 16'd11340;
          lut[9792] <= 16'd11467;
          lut[9793] <= 16'd11592;
          lut[9794] <= 16'd11716;
          lut[9795] <= 16'd11838;
          lut[9796] <= 16'd11959;
          lut[9797] <= 16'd12078;
          lut[9798] <= 16'd12195;
          lut[9799] <= 16'd12311;
          lut[9800] <= 16'd12425;
          lut[9801] <= 16'd12538;
          lut[9802] <= 16'd12650;
          lut[9803] <= 16'd12759;
          lut[9804] <= 16'd12868;
          lut[9805] <= 16'd12975;
          lut[9806] <= 16'd13081;
          lut[9807] <= 16'd13185;
          lut[9808] <= 16'd13288;
          lut[9809] <= 16'd13390;
          lut[9810] <= 16'd13490;
          lut[9811] <= 16'd13589;
          lut[9812] <= 16'd13686;
          lut[9813] <= 16'd13783;
          lut[9814] <= 16'd13878;
          lut[9815] <= 16'd13972;
          lut[9816] <= 16'd14065;
          lut[9817] <= 16'd14156;
          lut[9818] <= 16'd14246;
          lut[9819] <= 16'd14336;
          lut[9820] <= 16'd14424;
          lut[9821] <= 16'd14511;
          lut[9822] <= 16'd14596;
          lut[9823] <= 16'd14681;
          lut[9824] <= 16'd14765;
          lut[9825] <= 16'd14847;
          lut[9826] <= 16'd14929;
          lut[9827] <= 16'd15009;
          lut[9828] <= 16'd15088;
          lut[9829] <= 16'd15167;
          lut[9830] <= 16'd15244;
          lut[9831] <= 16'd15321;
          lut[9832] <= 16'd15396;
          lut[9833] <= 16'd15471;
          lut[9834] <= 16'd15545;
          lut[9835] <= 16'd15617;
          lut[9836] <= 16'd15689;
          lut[9837] <= 16'd15760;
          lut[9838] <= 16'd15830;
          lut[9839] <= 16'd15899;
          lut[9840] <= 16'd15968;
          lut[9841] <= 16'd16035;
          lut[9842] <= 16'd16102;
          lut[9843] <= 16'd16168;
          lut[9844] <= 16'd16233;
          lut[9845] <= 16'd16298;
          lut[9846] <= 16'd16361;
          lut[9847] <= 16'd16424;
          lut[9848] <= 16'd16486;
          lut[9849] <= 16'd16547;
          lut[9850] <= 16'd16608;
          lut[9851] <= 16'd16668;
          lut[9852] <= 16'd16727;
          lut[9853] <= 16'd16786;
          lut[9854] <= 16'd16844;
          lut[9855] <= 16'd16901;
          lut[9856] <= 0;
          lut[9857] <= 16'd213;
          lut[9858] <= 16'd425;
          lut[9859] <= 16'd638;
          lut[9860] <= 16'd850;
          lut[9861] <= 16'd1062;
          lut[9862] <= 16'd1274;
          lut[9863] <= 16'd1485;
          lut[9864] <= 16'd1696;
          lut[9865] <= 16'd1906;
          lut[9866] <= 16'd2116;
          lut[9867] <= 16'd2325;
          lut[9868] <= 16'd2533;
          lut[9869] <= 16'd2740;
          lut[9870] <= 16'd2947;
          lut[9871] <= 16'd3152;
          lut[9872] <= 16'd3357;
          lut[9873] <= 16'd3560;
          lut[9874] <= 16'd3762;
          lut[9875] <= 16'd3964;
          lut[9876] <= 16'd4164;
          lut[9877] <= 16'd4362;
          lut[9878] <= 16'd4560;
          lut[9879] <= 16'd4756;
          lut[9880] <= 16'd4950;
          lut[9881] <= 16'd5144;
          lut[9882] <= 16'd5335;
          lut[9883] <= 16'd5526;
          lut[9884] <= 16'd5714;
          lut[9885] <= 16'd5901;
          lut[9886] <= 16'd6087;
          lut[9887] <= 16'd6271;
          lut[9888] <= 16'd6453;
          lut[9889] <= 16'd6634;
          lut[9890] <= 16'd6813;
          lut[9891] <= 16'd6990;
          lut[9892] <= 16'd7165;
          lut[9893] <= 16'd7339;
          lut[9894] <= 16'd7511;
          lut[9895] <= 16'd7681;
          lut[9896] <= 16'd7850;
          lut[9897] <= 16'd8016;
          lut[9898] <= 16'd8181;
          lut[9899] <= 16'd8344;
          lut[9900] <= 16'd8506;
          lut[9901] <= 16'd8665;
          lut[9902] <= 16'd8823;
          lut[9903] <= 16'd8979;
          lut[9904] <= 16'd9133;
          lut[9905] <= 16'd9285;
          lut[9906] <= 16'd9436;
          lut[9907] <= 16'd9585;
          lut[9908] <= 16'd9732;
          lut[9909] <= 16'd9877;
          lut[9910] <= 16'd10020;
          lut[9911] <= 16'd10162;
          lut[9912] <= 16'd10302;
          lut[9913] <= 16'd10441;
          lut[9914] <= 16'd10577;
          lut[9915] <= 16'd10712;
          lut[9916] <= 16'd10845;
          lut[9917] <= 16'd10977;
          lut[9918] <= 16'd11107;
          lut[9919] <= 16'd11235;
          lut[9920] <= 16'd11362;
          lut[9921] <= 16'd11487;
          lut[9922] <= 16'd11610;
          lut[9923] <= 16'd11732;
          lut[9924] <= 16'd11852;
          lut[9925] <= 16'd11971;
          lut[9926] <= 16'd12088;
          lut[9927] <= 16'd12204;
          lut[9928] <= 16'd12318;
          lut[9929] <= 16'd12431;
          lut[9930] <= 16'd12542;
          lut[9931] <= 16'd12652;
          lut[9932] <= 16'd12761;
          lut[9933] <= 16'd12868;
          lut[9934] <= 16'd12974;
          lut[9935] <= 16'd13078;
          lut[9936] <= 16'd13181;
          lut[9937] <= 16'd13283;
          lut[9938] <= 16'd13383;
          lut[9939] <= 16'd13482;
          lut[9940] <= 16'd13580;
          lut[9941] <= 16'd13676;
          lut[9942] <= 16'd13772;
          lut[9943] <= 16'd13866;
          lut[9944] <= 16'd13959;
          lut[9945] <= 16'd14050;
          lut[9946] <= 16'd14141;
          lut[9947] <= 16'd14230;
          lut[9948] <= 16'd14318;
          lut[9949] <= 16'd14405;
          lut[9950] <= 16'd14491;
          lut[9951] <= 16'd14576;
          lut[9952] <= 16'd14660;
          lut[9953] <= 16'd14743;
          lut[9954] <= 16'd14825;
          lut[9955] <= 16'd14905;
          lut[9956] <= 16'd14985;
          lut[9957] <= 16'd15064;
          lut[9958] <= 16'd15142;
          lut[9959] <= 16'd15218;
          lut[9960] <= 16'd15294;
          lut[9961] <= 16'd15369;
          lut[9962] <= 16'd15443;
          lut[9963] <= 16'd15516;
          lut[9964] <= 16'd15588;
          lut[9965] <= 16'd15659;
          lut[9966] <= 16'd15730;
          lut[9967] <= 16'd15799;
          lut[9968] <= 16'd15868;
          lut[9969] <= 16'd15936;
          lut[9970] <= 16'd16003;
          lut[9971] <= 16'd16069;
          lut[9972] <= 16'd16135;
          lut[9973] <= 16'd16199;
          lut[9974] <= 16'd16263;
          lut[9975] <= 16'd16327;
          lut[9976] <= 16'd16389;
          lut[9977] <= 16'd16451;
          lut[9978] <= 16'd16512;
          lut[9979] <= 16'd16572;
          lut[9980] <= 16'd16631;
          lut[9981] <= 16'd16690;
          lut[9982] <= 16'd16748;
          lut[9983] <= 16'd16806;
          lut[9984] <= 0;
          lut[9985] <= 16'd210;
          lut[9986] <= 16'd420;
          lut[9987] <= 16'd630;
          lut[9988] <= 16'd839;
          lut[9989] <= 16'd1049;
          lut[9990] <= 16'd1258;
          lut[9991] <= 16'd1466;
          lut[9992] <= 16'd1675;
          lut[9993] <= 16'd1882;
          lut[9994] <= 16'd2089;
          lut[9995] <= 16'd2295;
          lut[9996] <= 16'd2501;
          lut[9997] <= 16'd2706;
          lut[9998] <= 16'd2910;
          lut[9999] <= 16'd3113;
          lut[10000] <= 16'd3315;
          lut[10001] <= 16'd3516;
          lut[10002] <= 16'd3716;
          lut[10003] <= 16'd3915;
          lut[10004] <= 16'd4112;
          lut[10005] <= 16'd4309;
          lut[10006] <= 16'd4504;
          lut[10007] <= 16'd4698;
          lut[10008] <= 16'd4891;
          lut[10009] <= 16'd5082;
          lut[10010] <= 16'd5272;
          lut[10011] <= 16'd5460;
          lut[10012] <= 16'd5647;
          lut[10013] <= 16'd5832;
          lut[10014] <= 16'd6016;
          lut[10015] <= 16'd6198;
          lut[10016] <= 16'd6379;
          lut[10017] <= 16'd6558;
          lut[10018] <= 16'd6735;
          lut[10019] <= 16'd6911;
          lut[10020] <= 16'd7085;
          lut[10021] <= 16'd7257;
          lut[10022] <= 16'd7428;
          lut[10023] <= 16'd7596;
          lut[10024] <= 16'd7764;
          lut[10025] <= 16'd7929;
          lut[10026] <= 16'd8093;
          lut[10027] <= 16'd8255;
          lut[10028] <= 16'd8415;
          lut[10029] <= 16'd8573;
          lut[10030] <= 16'd8730;
          lut[10031] <= 16'd8885;
          lut[10032] <= 16'd9038;
          lut[10033] <= 16'd9190;
          lut[10034] <= 16'd9340;
          lut[10035] <= 16'd9488;
          lut[10036] <= 16'd9634;
          lut[10037] <= 16'd9778;
          lut[10038] <= 16'd9921;
          lut[10039] <= 16'd10062;
          lut[10040] <= 16'd10202;
          lut[10041] <= 16'd10340;
          lut[10042] <= 16'd10476;
          lut[10043] <= 16'd10610;
          lut[10044] <= 16'd10743;
          lut[10045] <= 16'd10874;
          lut[10046] <= 16'd11004;
          lut[10047] <= 16'd11132;
          lut[10048] <= 16'd11258;
          lut[10049] <= 16'd11383;
          lut[10050] <= 16'd11506;
          lut[10051] <= 16'd11627;
          lut[10052] <= 16'd11748;
          lut[10053] <= 16'd11866;
          lut[10054] <= 16'd11983;
          lut[10055] <= 16'd12099;
          lut[10056] <= 16'd12213;
          lut[10057] <= 16'd12326;
          lut[10058] <= 16'd12437;
          lut[10059] <= 16'd12547;
          lut[10060] <= 16'd12655;
          lut[10061] <= 16'd12762;
          lut[10062] <= 16'd12868;
          lut[10063] <= 16'd12972;
          lut[10064] <= 16'd13075;
          lut[10065] <= 16'd13177;
          lut[10066] <= 16'd13277;
          lut[10067] <= 16'd13377;
          lut[10068] <= 16'd13475;
          lut[10069] <= 16'd13571;
          lut[10070] <= 16'd13667;
          lut[10071] <= 16'd13761;
          lut[10072] <= 16'd13854;
          lut[10073] <= 16'd13946;
          lut[10074] <= 16'd14036;
          lut[10075] <= 16'd14126;
          lut[10076] <= 16'd14214;
          lut[10077] <= 16'd14301;
          lut[10078] <= 16'd14388;
          lut[10079] <= 16'd14473;
          lut[10080] <= 16'd14557;
          lut[10081] <= 16'd14640;
          lut[10082] <= 16'd14722;
          lut[10083] <= 16'd14803;
          lut[10084] <= 16'd14883;
          lut[10085] <= 16'd14962;
          lut[10086] <= 16'd15040;
          lut[10087] <= 16'd15117;
          lut[10088] <= 16'd15193;
          lut[10089] <= 16'd15268;
          lut[10090] <= 16'd15342;
          lut[10091] <= 16'd15416;
          lut[10092] <= 16'd15488;
          lut[10093] <= 16'd15560;
          lut[10094] <= 16'd15630;
          lut[10095] <= 16'd15700;
          lut[10096] <= 16'd15769;
          lut[10097] <= 16'd15837;
          lut[10098] <= 16'd15905;
          lut[10099] <= 16'd15971;
          lut[10100] <= 16'd16037;
          lut[10101] <= 16'd16102;
          lut[10102] <= 16'd16166;
          lut[10103] <= 16'd16230;
          lut[10104] <= 16'd16293;
          lut[10105] <= 16'd16355;
          lut[10106] <= 16'd16416;
          lut[10107] <= 16'd16477;
          lut[10108] <= 16'd16536;
          lut[10109] <= 16'd16596;
          lut[10110] <= 16'd16654;
          lut[10111] <= 16'd16712;
          lut[10112] <= 0;
          lut[10113] <= 16'd207;
          lut[10114] <= 16'd415;
          lut[10115] <= 16'd622;
          lut[10116] <= 16'd829;
          lut[10117] <= 16'd1036;
          lut[10118] <= 16'd1242;
          lut[10119] <= 16'd1448;
          lut[10120] <= 16'd1654;
          lut[10121] <= 16'd1859;
          lut[10122] <= 16'd2063;
          lut[10123] <= 16'd2267;
          lut[10124] <= 16'd2470;
          lut[10125] <= 16'd2672;
          lut[10126] <= 16'd2874;
          lut[10127] <= 16'd3074;
          lut[10128] <= 16'd3274;
          lut[10129] <= 16'd3473;
          lut[10130] <= 16'd3670;
          lut[10131] <= 16'd3867;
          lut[10132] <= 16'd4062;
          lut[10133] <= 16'd4257;
          lut[10134] <= 16'd4450;
          lut[10135] <= 16'd4642;
          lut[10136] <= 16'd4832;
          lut[10137] <= 16'd5021;
          lut[10138] <= 16'd5209;
          lut[10139] <= 16'd5396;
          lut[10140] <= 16'd5581;
          lut[10141] <= 16'd5764;
          lut[10142] <= 16'd5946;
          lut[10143] <= 16'd6127;
          lut[10144] <= 16'd6306;
          lut[10145] <= 16'd6483;
          lut[10146] <= 16'd6659;
          lut[10147] <= 16'd6833;
          lut[10148] <= 16'd7005;
          lut[10149] <= 16'd7176;
          lut[10150] <= 16'd7346;
          lut[10151] <= 16'd7513;
          lut[10152] <= 16'd7679;
          lut[10153] <= 16'd7843;
          lut[10154] <= 16'd8006;
          lut[10155] <= 16'd8167;
          lut[10156] <= 16'd8326;
          lut[10157] <= 16'd8483;
          lut[10158] <= 16'd8639;
          lut[10159] <= 16'd8793;
          lut[10160] <= 16'd8945;
          lut[10161] <= 16'd9096;
          lut[10162] <= 16'd9245;
          lut[10163] <= 16'd9392;
          lut[10164] <= 16'd9538;
          lut[10165] <= 16'd9682;
          lut[10166] <= 16'd9824;
          lut[10167] <= 16'd9964;
          lut[10168] <= 16'd10103;
          lut[10169] <= 16'd10240;
          lut[10170] <= 16'd10376;
          lut[10171] <= 16'd10510;
          lut[10172] <= 16'd10642;
          lut[10173] <= 16'd10773;
          lut[10174] <= 16'd10902;
          lut[10175] <= 16'd11030;
          lut[10176] <= 16'd11156;
          lut[10177] <= 16'd11280;
          lut[10178] <= 16'd11403;
          lut[10179] <= 16'd11524;
          lut[10180] <= 16'd11644;
          lut[10181] <= 16'd11763;
          lut[10182] <= 16'd11880;
          lut[10183] <= 16'd11995;
          lut[10184] <= 16'd12109;
          lut[10185] <= 16'd12222;
          lut[10186] <= 16'd12333;
          lut[10187] <= 16'd12443;
          lut[10188] <= 16'd12551;
          lut[10189] <= 16'd12658;
          lut[10190] <= 16'd12764;
          lut[10191] <= 16'd12868;
          lut[10192] <= 16'd12971;
          lut[10193] <= 16'd13073;
          lut[10194] <= 16'd13173;
          lut[10195] <= 16'd13272;
          lut[10196] <= 16'd13370;
          lut[10197] <= 16'd13467;
          lut[10198] <= 16'd13563;
          lut[10199] <= 16'd13657;
          lut[10200] <= 16'd13750;
          lut[10201] <= 16'd13842;
          lut[10202] <= 16'd13933;
          lut[10203] <= 16'd14023;
          lut[10204] <= 16'd14111;
          lut[10205] <= 16'd14199;
          lut[10206] <= 16'd14285;
          lut[10207] <= 16'd14370;
          lut[10208] <= 16'd14455;
          lut[10209] <= 16'd14538;
          lut[10210] <= 16'd14620;
          lut[10211] <= 16'd14701;
          lut[10212] <= 16'd14781;
          lut[10213] <= 16'd14861;
          lut[10214] <= 16'd14939;
          lut[10215] <= 16'd15016;
          lut[10216] <= 16'd15092;
          lut[10217] <= 16'd15168;
          lut[10218] <= 16'd15242;
          lut[10219] <= 16'd15316;
          lut[10220] <= 16'd15389;
          lut[10221] <= 16'd15461;
          lut[10222] <= 16'd15532;
          lut[10223] <= 16'd15602;
          lut[10224] <= 16'd15671;
          lut[10225] <= 16'd15740;
          lut[10226] <= 16'd15807;
          lut[10227] <= 16'd15874;
          lut[10228] <= 16'd15940;
          lut[10229] <= 16'd16006;
          lut[10230] <= 16'd16070;
          lut[10231] <= 16'd16134;
          lut[10232] <= 16'd16197;
          lut[10233] <= 16'd16259;
          lut[10234] <= 16'd16321;
          lut[10235] <= 16'd16382;
          lut[10236] <= 16'd16442;
          lut[10237] <= 16'd16502;
          lut[10238] <= 16'd16560;
          lut[10239] <= 16'd16619;
          lut[10240] <= 0;
          lut[10241] <= 16'd205;
          lut[10242] <= 16'd410;
          lut[10243] <= 16'd614;
          lut[10244] <= 16'd819;
          lut[10245] <= 16'd1023;
          lut[10246] <= 16'd1227;
          lut[10247] <= 16'd1430;
          lut[10248] <= 16'd1633;
          lut[10249] <= 16'd1835;
          lut[10250] <= 16'd2037;
          lut[10251] <= 16'd2239;
          lut[10252] <= 16'd2439;
          lut[10253] <= 16'd2639;
          lut[10254] <= 16'd2838;
          lut[10255] <= 16'd3037;
          lut[10256] <= 16'd3234;
          lut[10257] <= 16'd3431;
          lut[10258] <= 16'd3626;
          lut[10259] <= 16'd3820;
          lut[10260] <= 16'd4014;
          lut[10261] <= 16'd4206;
          lut[10262] <= 16'd4397;
          lut[10263] <= 16'd4587;
          lut[10264] <= 16'd4775;
          lut[10265] <= 16'd4962;
          lut[10266] <= 16'd5148;
          lut[10267] <= 16'd5333;
          lut[10268] <= 16'd5516;
          lut[10269] <= 16'd5698;
          lut[10270] <= 16'd5878;
          lut[10271] <= 16'd6057;
          lut[10272] <= 16'd6234;
          lut[10273] <= 16'd6410;
          lut[10274] <= 16'd6584;
          lut[10275] <= 16'd6757;
          lut[10276] <= 16'd6928;
          lut[10277] <= 16'd7098;
          lut[10278] <= 16'd7265;
          lut[10279] <= 16'd7432;
          lut[10280] <= 16'd7596;
          lut[10281] <= 16'd7759;
          lut[10282] <= 16'd7921;
          lut[10283] <= 16'd8081;
          lut[10284] <= 16'd8239;
          lut[10285] <= 16'd8395;
          lut[10286] <= 16'd8550;
          lut[10287] <= 16'd8703;
          lut[10288] <= 16'd8854;
          lut[10289] <= 16'd9004;
          lut[10290] <= 16'd9152;
          lut[10291] <= 16'd9299;
          lut[10292] <= 16'd9443;
          lut[10293] <= 16'd9586;
          lut[10294] <= 16'd9728;
          lut[10295] <= 16'd9868;
          lut[10296] <= 16'd10006;
          lut[10297] <= 16'd10143;
          lut[10298] <= 16'd10278;
          lut[10299] <= 16'd10411;
          lut[10300] <= 16'd10543;
          lut[10301] <= 16'd10673;
          lut[10302] <= 16'd10802;
          lut[10303] <= 16'd10929;
          lut[10304] <= 16'd11055;
          lut[10305] <= 16'd11179;
          lut[10306] <= 16'd11302;
          lut[10307] <= 16'd11423;
          lut[10308] <= 16'd11542;
          lut[10309] <= 16'd11661;
          lut[10310] <= 16'd11777;
          lut[10311] <= 16'd11893;
          lut[10312] <= 16'd12006;
          lut[10313] <= 16'd12119;
          lut[10314] <= 16'd12230;
          lut[10315] <= 16'd12340;
          lut[10316] <= 16'd12448;
          lut[10317] <= 16'd12555;
          lut[10318] <= 16'd12661;
          lut[10319] <= 16'd12765;
          lut[10320] <= 16'd12868;
          lut[10321] <= 16'd12970;
          lut[10322] <= 16'd13070;
          lut[10323] <= 16'd13169;
          lut[10324] <= 16'd13267;
          lut[10325] <= 16'd13364;
          lut[10326] <= 16'd13460;
          lut[10327] <= 16'd13554;
          lut[10328] <= 16'd13648;
          lut[10329] <= 16'd13740;
          lut[10330] <= 16'd13831;
          lut[10331] <= 16'd13920;
          lut[10332] <= 16'd14009;
          lut[10333] <= 16'd14097;
          lut[10334] <= 16'd14183;
          lut[10335] <= 16'd14269;
          lut[10336] <= 16'd14353;
          lut[10337] <= 16'd14437;
          lut[10338] <= 16'd14519;
          lut[10339] <= 16'd14601;
          lut[10340] <= 16'd14681;
          lut[10341] <= 16'd14760;
          lut[10342] <= 16'd14839;
          lut[10343] <= 16'd14916;
          lut[10344] <= 16'd14993;
          lut[10345] <= 16'd15069;
          lut[10346] <= 16'd15143;
          lut[10347] <= 16'd15217;
          lut[10348] <= 16'd15290;
          lut[10349] <= 16'd15362;
          lut[10350] <= 16'd15434;
          lut[10351] <= 16'd15504;
          lut[10352] <= 16'd15574;
          lut[10353] <= 16'd15643;
          lut[10354] <= 16'd15711;
          lut[10355] <= 16'd15778;
          lut[10356] <= 16'd15844;
          lut[10357] <= 16'd15910;
          lut[10358] <= 16'd15975;
          lut[10359] <= 16'd16039;
          lut[10360] <= 16'd16102;
          lut[10361] <= 16'd16165;
          lut[10362] <= 16'd16227;
          lut[10363] <= 16'd16288;
          lut[10364] <= 16'd16348;
          lut[10365] <= 16'd16408;
          lut[10366] <= 16'd16467;
          lut[10367] <= 16'd16526;
          lut[10368] <= 0;
          lut[10369] <= 16'd202;
          lut[10370] <= 16'd404;
          lut[10371] <= 16'd607;
          lut[10372] <= 16'd808;
          lut[10373] <= 16'd1010;
          lut[10374] <= 16'd1211;
          lut[10375] <= 16'd1412;
          lut[10376] <= 16'd1613;
          lut[10377] <= 16'd1813;
          lut[10378] <= 16'd2013;
          lut[10379] <= 16'd2211;
          lut[10380] <= 16'd2410;
          lut[10381] <= 16'd2607;
          lut[10382] <= 16'd2804;
          lut[10383] <= 16'd3000;
          lut[10384] <= 16'd3195;
          lut[10385] <= 16'd3389;
          lut[10386] <= 16'd3583;
          lut[10387] <= 16'd3775;
          lut[10388] <= 16'd3966;
          lut[10389] <= 16'd4156;
          lut[10390] <= 16'd4345;
          lut[10391] <= 16'd4533;
          lut[10392] <= 16'd4720;
          lut[10393] <= 16'd4905;
          lut[10394] <= 16'd5089;
          lut[10395] <= 16'd5272;
          lut[10396] <= 16'd5453;
          lut[10397] <= 16'd5633;
          lut[10398] <= 16'd5811;
          lut[10399] <= 16'd5989;
          lut[10400] <= 16'd6164;
          lut[10401] <= 16'd6339;
          lut[10402] <= 16'd6511;
          lut[10403] <= 16'd6683;
          lut[10404] <= 16'd6852;
          lut[10405] <= 16'd7020;
          lut[10406] <= 16'd7187;
          lut[10407] <= 16'd7352;
          lut[10408] <= 16'd7515;
          lut[10409] <= 16'd7677;
          lut[10410] <= 16'd7837;
          lut[10411] <= 16'd7996;
          lut[10412] <= 16'd8153;
          lut[10413] <= 16'd8308;
          lut[10414] <= 16'd8462;
          lut[10415] <= 16'd8614;
          lut[10416] <= 16'd8765;
          lut[10417] <= 16'd8914;
          lut[10418] <= 16'd9061;
          lut[10419] <= 16'd9207;
          lut[10420] <= 16'd9351;
          lut[10421] <= 16'd9493;
          lut[10422] <= 16'd9634;
          lut[10423] <= 16'd9773;
          lut[10424] <= 16'd9911;
          lut[10425] <= 16'd10047;
          lut[10426] <= 16'd10181;
          lut[10427] <= 16'd10314;
          lut[10428] <= 16'd10446;
          lut[10429] <= 16'd10575;
          lut[10430] <= 16'd10704;
          lut[10431] <= 16'd10831;
          lut[10432] <= 16'd10956;
          lut[10433] <= 16'd11080;
          lut[10434] <= 16'd11202;
          lut[10435] <= 16'd11323;
          lut[10436] <= 16'd11442;
          lut[10437] <= 16'd11560;
          lut[10438] <= 16'd11677;
          lut[10439] <= 16'd11792;
          lut[10440] <= 16'd11905;
          lut[10441] <= 16'd12018;
          lut[10442] <= 16'd12129;
          lut[10443] <= 16'd12238;
          lut[10444] <= 16'd12346;
          lut[10445] <= 16'd12453;
          lut[10446] <= 16'd12559;
          lut[10447] <= 16'd12663;
          lut[10448] <= 16'd12766;
          lut[10449] <= 16'd12868;
          lut[10450] <= 16'd12968;
          lut[10451] <= 16'd13068;
          lut[10452] <= 16'd13166;
          lut[10453] <= 16'd13263;
          lut[10454] <= 16'd13358;
          lut[10455] <= 16'd13453;
          lut[10456] <= 16'd13546;
          lut[10457] <= 16'd13638;
          lut[10458] <= 16'd13729;
          lut[10459] <= 16'd13819;
          lut[10460] <= 16'd13908;
          lut[10461] <= 16'd13996;
          lut[10462] <= 16'd14083;
          lut[10463] <= 16'd14168;
          lut[10464] <= 16'd14253;
          lut[10465] <= 16'd14337;
          lut[10466] <= 16'd14419;
          lut[10467] <= 16'd14501;
          lut[10468] <= 16'd14582;
          lut[10469] <= 16'd14661;
          lut[10470] <= 16'd14740;
          lut[10471] <= 16'd14818;
          lut[10472] <= 16'd14894;
          lut[10473] <= 16'd14970;
          lut[10474] <= 16'd15045;
          lut[10475] <= 16'd15120;
          lut[10476] <= 16'd15193;
          lut[10477] <= 16'd15265;
          lut[10478] <= 16'd15337;
          lut[10479] <= 16'd15407;
          lut[10480] <= 16'd15477;
          lut[10481] <= 16'd15546;
          lut[10482] <= 16'd15615;
          lut[10483] <= 16'd15682;
          lut[10484] <= 16'd15749;
          lut[10485] <= 16'd15815;
          lut[10486] <= 16'd15880;
          lut[10487] <= 16'd15944;
          lut[10488] <= 16'd16008;
          lut[10489] <= 16'd16071;
          lut[10490] <= 16'd16133;
          lut[10491] <= 16'd16195;
          lut[10492] <= 16'd16255;
          lut[10493] <= 16'd16316;
          lut[10494] <= 16'd16375;
          lut[10495] <= 16'd16434;
          lut[10496] <= 0;
          lut[10497] <= 16'd200;
          lut[10498] <= 16'd400;
          lut[10499] <= 16'd599;
          lut[10500] <= 16'd799;
          lut[10501] <= 16'd998;
          lut[10502] <= 16'd1197;
          lut[10503] <= 16'd1395;
          lut[10504] <= 16'd1593;
          lut[10505] <= 16'd1791;
          lut[10506] <= 16'd1988;
          lut[10507] <= 16'd2185;
          lut[10508] <= 16'd2381;
          lut[10509] <= 16'd2576;
          lut[10510] <= 16'd2771;
          lut[10511] <= 16'd2964;
          lut[10512] <= 16'd3157;
          lut[10513] <= 16'd3349;
          lut[10514] <= 16'd3540;
          lut[10515] <= 16'd3730;
          lut[10516] <= 16'd3920;
          lut[10517] <= 16'd4108;
          lut[10518] <= 16'd4295;
          lut[10519] <= 16'd4480;
          lut[10520] <= 16'd4665;
          lut[10521] <= 16'd4848;
          lut[10522] <= 16'd5031;
          lut[10523] <= 16'd5212;
          lut[10524] <= 16'd5391;
          lut[10525] <= 16'd5569;
          lut[10526] <= 16'd5746;
          lut[10527] <= 16'd5922;
          lut[10528] <= 16'd6096;
          lut[10529] <= 16'd6269;
          lut[10530] <= 16'd6440;
          lut[10531] <= 16'd6610;
          lut[10532] <= 16'd6778;
          lut[10533] <= 16'd6945;
          lut[10534] <= 16'd7110;
          lut[10535] <= 16'd7274;
          lut[10536] <= 16'd7436;
          lut[10537] <= 16'd7596;
          lut[10538] <= 16'd7755;
          lut[10539] <= 16'd7913;
          lut[10540] <= 16'd8069;
          lut[10541] <= 16'd8223;
          lut[10542] <= 16'd8376;
          lut[10543] <= 16'd8527;
          lut[10544] <= 16'd8677;
          lut[10545] <= 16'd8825;
          lut[10546] <= 16'd8971;
          lut[10547] <= 16'd9116;
          lut[10548] <= 16'd9259;
          lut[10549] <= 16'd9401;
          lut[10550] <= 16'd9541;
          lut[10551] <= 16'd9680;
          lut[10552] <= 16'd9817;
          lut[10553] <= 16'd9952;
          lut[10554] <= 16'd10086;
          lut[10555] <= 16'd10219;
          lut[10556] <= 16'd10350;
          lut[10557] <= 16'd10479;
          lut[10558] <= 16'd10607;
          lut[10559] <= 16'd10733;
          lut[10560] <= 16'd10858;
          lut[10561] <= 16'd10982;
          lut[10562] <= 16'd11104;
          lut[10563] <= 16'd11224;
          lut[10564] <= 16'd11343;
          lut[10565] <= 16'd11461;
          lut[10566] <= 16'd11577;
          lut[10567] <= 16'd11692;
          lut[10568] <= 16'd11806;
          lut[10569] <= 16'd11918;
          lut[10570] <= 16'd12028;
          lut[10571] <= 16'd12138;
          lut[10572] <= 16'd12246;
          lut[10573] <= 16'd12353;
          lut[10574] <= 16'd12458;
          lut[10575] <= 16'd12563;
          lut[10576] <= 16'd12666;
          lut[10577] <= 16'd12767;
          lut[10578] <= 16'd12868;
          lut[10579] <= 16'd12967;
          lut[10580] <= 16'd13065;
          lut[10581] <= 16'd13162;
          lut[10582] <= 16'd13258;
          lut[10583] <= 16'd13353;
          lut[10584] <= 16'd13446;
          lut[10585] <= 16'd13538;
          lut[10586] <= 16'd13629;
          lut[10587] <= 16'd13720;
          lut[10588] <= 16'd13809;
          lut[10589] <= 16'd13896;
          lut[10590] <= 16'd13983;
          lut[10591] <= 16'd14069;
          lut[10592] <= 16'd14154;
          lut[10593] <= 16'd14238;
          lut[10594] <= 16'd14321;
          lut[10595] <= 16'd14402;
          lut[10596] <= 16'd14483;
          lut[10597] <= 16'd14563;
          lut[10598] <= 16'd14642;
          lut[10599] <= 16'd14720;
          lut[10600] <= 16'd14797;
          lut[10601] <= 16'd14873;
          lut[10602] <= 16'd14948;
          lut[10603] <= 16'd15023;
          lut[10604] <= 16'd15096;
          lut[10605] <= 16'd15169;
          lut[10606] <= 16'd15241;
          lut[10607] <= 16'd15312;
          lut[10608] <= 16'd15382;
          lut[10609] <= 16'd15451;
          lut[10610] <= 16'd15520;
          lut[10611] <= 16'd15587;
          lut[10612] <= 16'd15654;
          lut[10613] <= 16'd15720;
          lut[10614] <= 16'd15786;
          lut[10615] <= 16'd15851;
          lut[10616] <= 16'd15914;
          lut[10617] <= 16'd15978;
          lut[10618] <= 16'd16040;
          lut[10619] <= 16'd16102;
          lut[10620] <= 16'd16163;
          lut[10621] <= 16'd16224;
          lut[10622] <= 16'd16283;
          lut[10623] <= 16'd16343;
          lut[10624] <= 0;
          lut[10625] <= 16'd197;
          lut[10626] <= 16'd395;
          lut[10627] <= 16'd592;
          lut[10628] <= 16'd789;
          lut[10629] <= 16'd986;
          lut[10630] <= 16'd1182;
          lut[10631] <= 16'd1379;
          lut[10632] <= 16'd1574;
          lut[10633] <= 16'd1770;
          lut[10634] <= 16'd1965;
          lut[10635] <= 16'd2159;
          lut[10636] <= 16'd2352;
          lut[10637] <= 16'd2545;
          lut[10638] <= 16'd2738;
          lut[10639] <= 16'd2929;
          lut[10640] <= 16'd3120;
          lut[10641] <= 16'd3310;
          lut[10642] <= 16'd3499;
          lut[10643] <= 16'd3687;
          lut[10644] <= 16'd3874;
          lut[10645] <= 16'd4060;
          lut[10646] <= 16'd4245;
          lut[10647] <= 16'd4429;
          lut[10648] <= 16'd4612;
          lut[10649] <= 16'd4793;
          lut[10650] <= 16'd4974;
          lut[10651] <= 16'd5153;
          lut[10652] <= 16'd5331;
          lut[10653] <= 16'd5507;
          lut[10654] <= 16'd5683;
          lut[10655] <= 16'd5856;
          lut[10656] <= 16'd6029;
          lut[10657] <= 16'd6200;
          lut[10658] <= 16'd6370;
          lut[10659] <= 16'd6538;
          lut[10660] <= 16'd6705;
          lut[10661] <= 16'd6870;
          lut[10662] <= 16'd7034;
          lut[10663] <= 16'd7197;
          lut[10664] <= 16'd7358;
          lut[10665] <= 16'd7517;
          lut[10666] <= 16'd7675;
          lut[10667] <= 16'd7832;
          lut[10668] <= 16'd7986;
          lut[10669] <= 16'd8140;
          lut[10670] <= 16'd8292;
          lut[10671] <= 16'd8442;
          lut[10672] <= 16'd8590;
          lut[10673] <= 16'd8738;
          lut[10674] <= 16'd8883;
          lut[10675] <= 16'd9027;
          lut[10676] <= 16'd9170;
          lut[10677] <= 16'd9311;
          lut[10678] <= 16'd9450;
          lut[10679] <= 16'd9588;
          lut[10680] <= 16'd9725;
          lut[10681] <= 16'd9859;
          lut[10682] <= 16'd9993;
          lut[10683] <= 16'd10125;
          lut[10684] <= 16'd10255;
          lut[10685] <= 16'd10384;
          lut[10686] <= 16'd10511;
          lut[10687] <= 16'd10637;
          lut[10688] <= 16'd10762;
          lut[10689] <= 16'd10885;
          lut[10690] <= 16'd11007;
          lut[10691] <= 16'd11127;
          lut[10692] <= 16'd11246;
          lut[10693] <= 16'd11363;
          lut[10694] <= 16'd11479;
          lut[10695] <= 16'd11594;
          lut[10696] <= 16'd11707;
          lut[10697] <= 16'd11819;
          lut[10698] <= 16'd11930;
          lut[10699] <= 16'd12039;
          lut[10700] <= 16'd12147;
          lut[10701] <= 16'd12254;
          lut[10702] <= 16'd12359;
          lut[10703] <= 16'd12464;
          lut[10704] <= 16'd12566;
          lut[10705] <= 16'd12668;
          lut[10706] <= 16'd12769;
          lut[10707] <= 16'd12868;
          lut[10708] <= 16'd12966;
          lut[10709] <= 16'd13063;
          lut[10710] <= 16'd13159;
          lut[10711] <= 16'd13253;
          lut[10712] <= 16'd13347;
          lut[10713] <= 16'd13439;
          lut[10714] <= 16'd13531;
          lut[10715] <= 16'd13621;
          lut[10716] <= 16'd13710;
          lut[10717] <= 16'd13798;
          lut[10718] <= 16'd13885;
          lut[10719] <= 16'd13971;
          lut[10720] <= 16'd14056;
          lut[10721] <= 16'd14140;
          lut[10722] <= 16'd14223;
          lut[10723] <= 16'd14305;
          lut[10724] <= 16'd14386;
          lut[10725] <= 16'd14466;
          lut[10726] <= 16'd14545;
          lut[10727] <= 16'd14623;
          lut[10728] <= 16'd14700;
          lut[10729] <= 16'd14777;
          lut[10730] <= 16'd14852;
          lut[10731] <= 16'd14927;
          lut[10732] <= 16'd15000;
          lut[10733] <= 16'd15073;
          lut[10734] <= 16'd15145;
          lut[10735] <= 16'd15216;
          lut[10736] <= 16'd15287;
          lut[10737] <= 16'd15356;
          lut[10738] <= 16'd15425;
          lut[10739] <= 16'd15493;
          lut[10740] <= 16'd15560;
          lut[10741] <= 16'd15627;
          lut[10742] <= 16'd15693;
          lut[10743] <= 16'd15758;
          lut[10744] <= 16'd15822;
          lut[10745] <= 16'd15885;
          lut[10746] <= 16'd15948;
          lut[10747] <= 16'd16010;
          lut[10748] <= 16'd16072;
          lut[10749] <= 16'd16132;
          lut[10750] <= 16'd16192;
          lut[10751] <= 16'd16252;
          lut[10752] <= 0;
          lut[10753] <= 16'd195;
          lut[10754] <= 16'd390;
          lut[10755] <= 16'd585;
          lut[10756] <= 16'd780;
          lut[10757] <= 16'd974;
          lut[10758] <= 16'd1168;
          lut[10759] <= 16'd1362;
          lut[10760] <= 16'd1556;
          lut[10761] <= 16'd1749;
          lut[10762] <= 16'd1941;
          lut[10763] <= 16'd2133;
          lut[10764] <= 16'd2325;
          lut[10765] <= 16'd2516;
          lut[10766] <= 16'd2706;
          lut[10767] <= 16'd2895;
          lut[10768] <= 16'd3084;
          lut[10769] <= 16'd3272;
          lut[10770] <= 16'd3459;
          lut[10771] <= 16'd3645;
          lut[10772] <= 16'd3830;
          lut[10773] <= 16'd4014;
          lut[10774] <= 16'd4197;
          lut[10775] <= 16'd4379;
          lut[10776] <= 16'd4560;
          lut[10777] <= 16'd4739;
          lut[10778] <= 16'd4918;
          lut[10779] <= 16'd5095;
          lut[10780] <= 16'd5272;
          lut[10781] <= 16'd5446;
          lut[10782] <= 16'd5620;
          lut[10783] <= 16'd5792;
          lut[10784] <= 16'd5963;
          lut[10785] <= 16'd6133;
          lut[10786] <= 16'd6301;
          lut[10787] <= 16'd6468;
          lut[10788] <= 16'd6634;
          lut[10789] <= 16'd6798;
          lut[10790] <= 16'd6960;
          lut[10791] <= 16'd7122;
          lut[10792] <= 16'd7281;
          lut[10793] <= 16'd7440;
          lut[10794] <= 16'd7596;
          lut[10795] <= 16'd7752;
          lut[10796] <= 16'd7905;
          lut[10797] <= 16'd8058;
          lut[10798] <= 16'd8209;
          lut[10799] <= 16'd8358;
          lut[10800] <= 16'd8506;
          lut[10801] <= 16'd8652;
          lut[10802] <= 16'd8797;
          lut[10803] <= 16'd8940;
          lut[10804] <= 16'd9082;
          lut[10805] <= 16'd9222;
          lut[10806] <= 16'd9361;
          lut[10807] <= 16'd9498;
          lut[10808] <= 16'd9634;
          lut[10809] <= 16'd9768;
          lut[10810] <= 16'd9901;
          lut[10811] <= 16'd10032;
          lut[10812] <= 16'd10162;
          lut[10813] <= 16'd10291;
          lut[10814] <= 16'd10418;
          lut[10815] <= 16'd10543;
          lut[10816] <= 16'd10667;
          lut[10817] <= 16'd10790;
          lut[10818] <= 16'd10911;
          lut[10819] <= 16'd11031;
          lut[10820] <= 16'd11150;
          lut[10821] <= 16'd11267;
          lut[10822] <= 16'd11383;
          lut[10823] <= 16'd11497;
          lut[10824] <= 16'd11610;
          lut[10825] <= 16'd11722;
          lut[10826] <= 16'd11832;
          lut[10827] <= 16'd11942;
          lut[10828] <= 16'd12049;
          lut[10829] <= 16'd12156;
          lut[10830] <= 16'd12261;
          lut[10831] <= 16'd12366;
          lut[10832] <= 16'd12468;
          lut[10833] <= 16'd12570;
          lut[10834] <= 16'd12671;
          lut[10835] <= 16'd12770;
          lut[10836] <= 16'd12868;
          lut[10837] <= 16'd12965;
          lut[10838] <= 16'd13061;
          lut[10839] <= 16'd13155;
          lut[10840] <= 16'd13249;
          lut[10841] <= 16'd13341;
          lut[10842] <= 16'd13433;
          lut[10843] <= 16'd13523;
          lut[10844] <= 16'd13612;
          lut[10845] <= 16'd13700;
          lut[10846] <= 16'd13787;
          lut[10847] <= 16'd13874;
          lut[10848] <= 16'd13959;
          lut[10849] <= 16'd14043;
          lut[10850] <= 16'd14126;
          lut[10851] <= 16'd14208;
          lut[10852] <= 16'd14289;
          lut[10853] <= 16'd14369;
          lut[10854] <= 16'd14449;
          lut[10855] <= 16'd14527;
          lut[10856] <= 16'd14604;
          lut[10857] <= 16'd14681;
          lut[10858] <= 16'd14757;
          lut[10859] <= 16'd14831;
          lut[10860] <= 16'd14905;
          lut[10861] <= 16'd14978;
          lut[10862] <= 16'd15051;
          lut[10863] <= 16'd15122;
          lut[10864] <= 16'd15193;
          lut[10865] <= 16'd15263;
          lut[10866] <= 16'd15332;
          lut[10867] <= 16'd15400;
          lut[10868] <= 16'd15467;
          lut[10869] <= 16'd15534;
          lut[10870] <= 16'd15600;
          lut[10871] <= 16'd15665;
          lut[10872] <= 16'd15730;
          lut[10873] <= 16'd15794;
          lut[10874] <= 16'd15857;
          lut[10875] <= 16'd15919;
          lut[10876] <= 16'd15981;
          lut[10877] <= 16'd16042;
          lut[10878] <= 16'd16102;
          lut[10879] <= 16'd16162;
          lut[10880] <= 0;
          lut[10881] <= 16'd193;
          lut[10882] <= 16'd385;
          lut[10883] <= 16'd578;
          lut[10884] <= 16'd770;
          lut[10885] <= 16'd963;
          lut[10886] <= 16'd1155;
          lut[10887] <= 16'd1346;
          lut[10888] <= 16'd1537;
          lut[10889] <= 16'd1728;
          lut[10890] <= 16'd1919;
          lut[10891] <= 16'd2109;
          lut[10892] <= 16'd2298;
          lut[10893] <= 16'd2487;
          lut[10894] <= 16'd2675;
          lut[10895] <= 16'd2862;
          lut[10896] <= 16'd3048;
          lut[10897] <= 16'd3234;
          lut[10898] <= 16'd3419;
          lut[10899] <= 16'd3603;
          lut[10900] <= 16'd3786;
          lut[10901] <= 16'd3968;
          lut[10902] <= 16'd4150;
          lut[10903] <= 16'd4330;
          lut[10904] <= 16'd4509;
          lut[10905] <= 16'd4687;
          lut[10906] <= 16'd4864;
          lut[10907] <= 16'd5039;
          lut[10908] <= 16'd5214;
          lut[10909] <= 16'd5387;
          lut[10910] <= 16'd5559;
          lut[10911] <= 16'd5730;
          lut[10912] <= 16'd5899;
          lut[10913] <= 16'd6067;
          lut[10914] <= 16'd6234;
          lut[10915] <= 16'd6400;
          lut[10916] <= 16'd6564;
          lut[10917] <= 16'd6727;
          lut[10918] <= 16'd6888;
          lut[10919] <= 16'd7048;
          lut[10920] <= 16'd7206;
          lut[10921] <= 16'd7363;
          lut[10922] <= 16'd7519;
          lut[10923] <= 16'd7673;
          lut[10924] <= 16'd7826;
          lut[10925] <= 16'd7977;
          lut[10926] <= 16'd8127;
          lut[10927] <= 16'd8276;
          lut[10928] <= 16'd8422;
          lut[10929] <= 16'd8568;
          lut[10930] <= 16'd8712;
          lut[10931] <= 16'd8854;
          lut[10932] <= 16'd8995;
          lut[10933] <= 16'd9135;
          lut[10934] <= 16'd9273;
          lut[10935] <= 16'd9409;
          lut[10936] <= 16'd9545;
          lut[10937] <= 16'd9678;
          lut[10938] <= 16'd9810;
          lut[10939] <= 16'd9941;
          lut[10940] <= 16'd10071;
          lut[10941] <= 16'd10199;
          lut[10942] <= 16'd10325;
          lut[10943] <= 16'd10450;
          lut[10944] <= 16'd10574;
          lut[10945] <= 16'd10696;
          lut[10946] <= 16'd10817;
          lut[10947] <= 16'd10937;
          lut[10948] <= 16'd11055;
          lut[10949] <= 16'd11172;
          lut[10950] <= 16'd11287;
          lut[10951] <= 16'd11402;
          lut[10952] <= 16'd11514;
          lut[10953] <= 16'd11626;
          lut[10954] <= 16'd11736;
          lut[10955] <= 16'd11845;
          lut[10956] <= 16'd11953;
          lut[10957] <= 16'd12060;
          lut[10958] <= 16'd12165;
          lut[10959] <= 16'd12269;
          lut[10960] <= 16'd12372;
          lut[10961] <= 16'd12473;
          lut[10962] <= 16'd12574;
          lut[10963] <= 16'd12673;
          lut[10964] <= 16'd12771;
          lut[10965] <= 16'd12868;
          lut[10966] <= 16'd12964;
          lut[10967] <= 16'd13058;
          lut[10968] <= 16'd13152;
          lut[10969] <= 16'd13245;
          lut[10970] <= 16'd13336;
          lut[10971] <= 16'd13426;
          lut[10972] <= 16'd13516;
          lut[10973] <= 16'd13604;
          lut[10974] <= 16'd13691;
          lut[10975] <= 16'd13777;
          lut[10976] <= 16'd13862;
          lut[10977] <= 16'd13947;
          lut[10978] <= 16'd14030;
          lut[10979] <= 16'd14112;
          lut[10980] <= 16'd14193;
          lut[10981] <= 16'd14274;
          lut[10982] <= 16'd14353;
          lut[10983] <= 16'd14432;
          lut[10984] <= 16'd14510;
          lut[10985] <= 16'd14586;
          lut[10986] <= 16'd14662;
          lut[10987] <= 16'd14737;
          lut[10988] <= 16'd14811;
          lut[10989] <= 16'd14885;
          lut[10990] <= 16'd14957;
          lut[10991] <= 16'd15029;
          lut[10992] <= 16'd15100;
          lut[10993] <= 16'd15170;
          lut[10994] <= 16'd15239;
          lut[10995] <= 16'd15307;
          lut[10996] <= 16'd15375;
          lut[10997] <= 16'd15442;
          lut[10998] <= 16'd15508;
          lut[10999] <= 16'd15574;
          lut[11000] <= 16'd15639;
          lut[11001] <= 16'd15703;
          lut[11002] <= 16'd15766;
          lut[11003] <= 16'd15829;
          lut[11004] <= 16'd15891;
          lut[11005] <= 16'd15952;
          lut[11006] <= 16'd16012;
          lut[11007] <= 16'd16072;
          lut[11008] <= 0;
          lut[11009] <= 16'd191;
          lut[11010] <= 16'd381;
          lut[11011] <= 16'd571;
          lut[11012] <= 16'd761;
          lut[11013] <= 16'd951;
          lut[11014] <= 16'd1141;
          lut[11015] <= 16'd1331;
          lut[11016] <= 16'd1520;
          lut[11017] <= 16'd1708;
          lut[11018] <= 16'd1897;
          lut[11019] <= 16'd2084;
          lut[11020] <= 16'd2271;
          lut[11021] <= 16'd2458;
          lut[11022] <= 16'd2644;
          lut[11023] <= 16'd2829;
          lut[11024] <= 16'd3014;
          lut[11025] <= 16'd3197;
          lut[11026] <= 16'd3380;
          lut[11027] <= 16'd3562;
          lut[11028] <= 16'd3744;
          lut[11029] <= 16'd3924;
          lut[11030] <= 16'd4103;
          lut[11031] <= 16'd4282;
          lut[11032] <= 16'd4459;
          lut[11033] <= 16'd4635;
          lut[11034] <= 16'd4810;
          lut[11035] <= 16'd4984;
          lut[11036] <= 16'd5157;
          lut[11037] <= 16'd5329;
          lut[11038] <= 16'd5499;
          lut[11039] <= 16'd5668;
          lut[11040] <= 16'd5836;
          lut[11041] <= 16'd6003;
          lut[11042] <= 16'd6168;
          lut[11043] <= 16'd6333;
          lut[11044] <= 16'd6495;
          lut[11045] <= 16'd6657;
          lut[11046] <= 16'd6817;
          lut[11047] <= 16'd6976;
          lut[11048] <= 16'd7133;
          lut[11049] <= 16'd7289;
          lut[11050] <= 16'd7443;
          lut[11051] <= 16'd7596;
          lut[11052] <= 16'd7748;
          lut[11053] <= 16'd7898;
          lut[11054] <= 16'd8047;
          lut[11055] <= 16'd8195;
          lut[11056] <= 16'd8341;
          lut[11057] <= 16'd8485;
          lut[11058] <= 16'd8628;
          lut[11059] <= 16'd8770;
          lut[11060] <= 16'd8910;
          lut[11061] <= 16'd9049;
          lut[11062] <= 16'd9186;
          lut[11063] <= 16'd9322;
          lut[11064] <= 16'd9457;
          lut[11065] <= 16'd9590;
          lut[11066] <= 16'd9721;
          lut[11067] <= 16'd9852;
          lut[11068] <= 16'd9981;
          lut[11069] <= 16'd10108;
          lut[11070] <= 16'd10234;
          lut[11071] <= 16'd10359;
          lut[11072] <= 16'd10482;
          lut[11073] <= 16'd10604;
          lut[11074] <= 16'd10724;
          lut[11075] <= 16'd10844;
          lut[11076] <= 16'd10962;
          lut[11077] <= 16'd11078;
          lut[11078] <= 16'd11193;
          lut[11079] <= 16'd11307;
          lut[11080] <= 16'd11420;
          lut[11081] <= 16'd11531;
          lut[11082] <= 16'd11641;
          lut[11083] <= 16'd11750;
          lut[11084] <= 16'd11858;
          lut[11085] <= 16'd11964;
          lut[11086] <= 16'd12069;
          lut[11087] <= 16'd12173;
          lut[11088] <= 16'd12276;
          lut[11089] <= 16'd12378;
          lut[11090] <= 16'd12478;
          lut[11091] <= 16'd12577;
          lut[11092] <= 16'd12675;
          lut[11093] <= 16'd12772;
          lut[11094] <= 16'd12868;
          lut[11095] <= 16'd12963;
          lut[11096] <= 16'd13056;
          lut[11097] <= 16'd13149;
          lut[11098] <= 16'd13240;
          lut[11099] <= 16'd13331;
          lut[11100] <= 16'd13420;
          lut[11101] <= 16'd13508;
          lut[11102] <= 16'd13596;
          lut[11103] <= 16'd13682;
          lut[11104] <= 16'd13767;
          lut[11105] <= 16'd13852;
          lut[11106] <= 16'd13935;
          lut[11107] <= 16'd14017;
          lut[11108] <= 16'd14099;
          lut[11109] <= 16'd14179;
          lut[11110] <= 16'd14259;
          lut[11111] <= 16'd14338;
          lut[11112] <= 16'd14416;
          lut[11113] <= 16'd14492;
          lut[11114] <= 16'd14568;
          lut[11115] <= 16'd14644;
          lut[11116] <= 16'd14718;
          lut[11117] <= 16'd14792;
          lut[11118] <= 16'd14864;
          lut[11119] <= 16'd14936;
          lut[11120] <= 16'd15007;
          lut[11121] <= 16'd15077;
          lut[11122] <= 16'd15147;
          lut[11123] <= 16'd15216;
          lut[11124] <= 16'd15284;
          lut[11125] <= 16'd15351;
          lut[11126] <= 16'd15417;
          lut[11127] <= 16'd15483;
          lut[11128] <= 16'd15548;
          lut[11129] <= 16'd15612;
          lut[11130] <= 16'd15676;
          lut[11131] <= 16'd15739;
          lut[11132] <= 16'd15801;
          lut[11133] <= 16'd15862;
          lut[11134] <= 16'd15923;
          lut[11135] <= 16'd15984;
          lut[11136] <= 0;
          lut[11137] <= 16'd188;
          lut[11138] <= 16'd377;
          lut[11139] <= 16'd565;
          lut[11140] <= 16'd753;
          lut[11141] <= 16'd941;
          lut[11142] <= 16'd1128;
          lut[11143] <= 16'd1315;
          lut[11144] <= 16'd1502;
          lut[11145] <= 16'd1689;
          lut[11146] <= 16'd1875;
          lut[11147] <= 16'd2061;
          lut[11148] <= 16'd2246;
          lut[11149] <= 16'd2430;
          lut[11150] <= 16'd2614;
          lut[11151] <= 16'd2797;
          lut[11152] <= 16'd2980;
          lut[11153] <= 16'd3162;
          lut[11154] <= 16'd3343;
          lut[11155] <= 16'd3523;
          lut[11156] <= 16'd3702;
          lut[11157] <= 16'd3881;
          lut[11158] <= 16'd4058;
          lut[11159] <= 16'd4235;
          lut[11160] <= 16'd4410;
          lut[11161] <= 16'd4585;
          lut[11162] <= 16'd4758;
          lut[11163] <= 16'd4930;
          lut[11164] <= 16'd5101;
          lut[11165] <= 16'd5272;
          lut[11166] <= 16'd5440;
          lut[11167] <= 16'd5608;
          lut[11168] <= 16'd5775;
          lut[11169] <= 16'd5940;
          lut[11170] <= 16'd6104;
          lut[11171] <= 16'd6267;
          lut[11172] <= 16'd6428;
          lut[11173] <= 16'd6588;
          lut[11174] <= 16'd6747;
          lut[11175] <= 16'd6905;
          lut[11176] <= 16'd7061;
          lut[11177] <= 16'd7215;
          lut[11178] <= 16'd7369;
          lut[11179] <= 16'd7521;
          lut[11180] <= 16'd7672;
          lut[11181] <= 16'd7821;
          lut[11182] <= 16'd7969;
          lut[11183] <= 16'd8115;
          lut[11184] <= 16'd8260;
          lut[11185] <= 16'd8404;
          lut[11186] <= 16'd8546;
          lut[11187] <= 16'd8687;
          lut[11188] <= 16'd8827;
          lut[11189] <= 16'd8965;
          lut[11190] <= 16'd9101;
          lut[11191] <= 16'd9236;
          lut[11192] <= 16'd9370;
          lut[11193] <= 16'd9503;
          lut[11194] <= 16'd9634;
          lut[11195] <= 16'd9764;
          lut[11196] <= 16'd9892;
          lut[11197] <= 16'd10019;
          lut[11198] <= 16'd10144;
          lut[11199] <= 16'd10269;
          lut[11200] <= 16'd10391;
          lut[11201] <= 16'd10513;
          lut[11202] <= 16'd10633;
          lut[11203] <= 16'd10752;
          lut[11204] <= 16'd10870;
          lut[11205] <= 16'd10986;
          lut[11206] <= 16'd11101;
          lut[11207] <= 16'd11214;
          lut[11208] <= 16'd11327;
          lut[11209] <= 16'd11438;
          lut[11210] <= 16'd11548;
          lut[11211] <= 16'd11657;
          lut[11212] <= 16'd11764;
          lut[11213] <= 16'd11870;
          lut[11214] <= 16'd11975;
          lut[11215] <= 16'd12079;
          lut[11216] <= 16'd12182;
          lut[11217] <= 16'd12283;
          lut[11218] <= 16'd12383;
          lut[11219] <= 16'd12483;
          lut[11220] <= 16'd12581;
          lut[11221] <= 16'd12677;
          lut[11222] <= 16'd12773;
          lut[11223] <= 16'd12868;
          lut[11224] <= 16'd12962;
          lut[11225] <= 16'd13054;
          lut[11226] <= 16'd13146;
          lut[11227] <= 16'd13236;
          lut[11228] <= 16'd13325;
          lut[11229] <= 16'd13414;
          lut[11230] <= 16'd13501;
          lut[11231] <= 16'd13588;
          lut[11232] <= 16'd13673;
          lut[11233] <= 16'd13758;
          lut[11234] <= 16'd13841;
          lut[11235] <= 16'd13924;
          lut[11236] <= 16'd14005;
          lut[11237] <= 16'd14086;
          lut[11238] <= 16'd14166;
          lut[11239] <= 16'd14244;
          lut[11240] <= 16'd14322;
          lut[11241] <= 16'd14399;
          lut[11242] <= 16'd14476;
          lut[11243] <= 16'd14551;
          lut[11244] <= 16'd14626;
          lut[11245] <= 16'd14699;
          lut[11246] <= 16'd14772;
          lut[11247] <= 16'd14844;
          lut[11248] <= 16'd14916;
          lut[11249] <= 16'd14986;
          lut[11250] <= 16'd15056;
          lut[11251] <= 16'd15125;
          lut[11252] <= 16'd15193;
          lut[11253] <= 16'd15260;
          lut[11254] <= 16'd15327;
          lut[11255] <= 16'd15393;
          lut[11256] <= 16'd15458;
          lut[11257] <= 16'd15523;
          lut[11258] <= 16'd15586;
          lut[11259] <= 16'd15650;
          lut[11260] <= 16'd15712;
          lut[11261] <= 16'd15774;
          lut[11262] <= 16'd15835;
          lut[11263] <= 16'd15895;
          lut[11264] <= 0;
          lut[11265] <= 16'd186;
          lut[11266] <= 16'd372;
          lut[11267] <= 16'd558;
          lut[11268] <= 16'd744;
          lut[11269] <= 16'd930;
          lut[11270] <= 16'd1115;
          lut[11271] <= 16'd1301;
          lut[11272] <= 16'd1485;
          lut[11273] <= 16'd1670;
          lut[11274] <= 16'd1854;
          lut[11275] <= 16'd2037;
          lut[11276] <= 16'd2220;
          lut[11277] <= 16'd2403;
          lut[11278] <= 16'd2585;
          lut[11279] <= 16'd2766;
          lut[11280] <= 16'd2947;
          lut[11281] <= 16'd3127;
          lut[11282] <= 16'd3306;
          lut[11283] <= 16'd3484;
          lut[11284] <= 16'd3661;
          lut[11285] <= 16'd3838;
          lut[11286] <= 16'd4014;
          lut[11287] <= 16'd4188;
          lut[11288] <= 16'd4362;
          lut[11289] <= 16'd4535;
          lut[11290] <= 16'd4707;
          lut[11291] <= 16'd4878;
          lut[11292] <= 16'd5047;
          lut[11293] <= 16'd5216;
          lut[11294] <= 16'd5383;
          lut[11295] <= 16'd5549;
          lut[11296] <= 16'd5714;
          lut[11297] <= 16'd5878;
          lut[11298] <= 16'd6041;
          lut[11299] <= 16'd6202;
          lut[11300] <= 16'd6362;
          lut[11301] <= 16'd6521;
          lut[11302] <= 16'd6679;
          lut[11303] <= 16'd6835;
          lut[11304] <= 16'd6990;
          lut[11305] <= 16'd7144;
          lut[11306] <= 16'd7296;
          lut[11307] <= 16'd7447;
          lut[11308] <= 16'd7596;
          lut[11309] <= 16'd7745;
          lut[11310] <= 16'd7892;
          lut[11311] <= 16'd8037;
          lut[11312] <= 16'd8181;
          lut[11313] <= 16'd8324;
          lut[11314] <= 16'd8466;
          lut[11315] <= 16'd8606;
          lut[11316] <= 16'd8744;
          lut[11317] <= 16'd8882;
          lut[11318] <= 16'd9018;
          lut[11319] <= 16'd9152;
          lut[11320] <= 16'd9285;
          lut[11321] <= 16'd9417;
          lut[11322] <= 16'd9548;
          lut[11323] <= 16'd9677;
          lut[11324] <= 16'd9804;
          lut[11325] <= 16'd9931;
          lut[11326] <= 16'd10056;
          lut[11327] <= 16'd10180;
          lut[11328] <= 16'd10302;
          lut[11329] <= 16'd10423;
          lut[11330] <= 16'd10543;
          lut[11331] <= 16'd10662;
          lut[11332] <= 16'd10779;
          lut[11333] <= 16'd10895;
          lut[11334] <= 16'd11009;
          lut[11335] <= 16'd11123;
          lut[11336] <= 16'd11235;
          lut[11337] <= 16'd11346;
          lut[11338] <= 16'd11456;
          lut[11339] <= 16'd11564;
          lut[11340] <= 16'd11671;
          lut[11341] <= 16'd11777;
          lut[11342] <= 16'd11882;
          lut[11343] <= 16'd11986;
          lut[11344] <= 16'd12088;
          lut[11345] <= 16'd12190;
          lut[11346] <= 16'd12290;
          lut[11347] <= 16'd12389;
          lut[11348] <= 16'd12487;
          lut[11349] <= 16'd12584;
          lut[11350] <= 16'd12680;
          lut[11351] <= 16'd12774;
          lut[11352] <= 16'd12868;
          lut[11353] <= 16'd12961;
          lut[11354] <= 16'd13052;
          lut[11355] <= 16'd13143;
          lut[11356] <= 16'd13232;
          lut[11357] <= 16'd13320;
          lut[11358] <= 16'd13408;
          lut[11359] <= 16'd13494;
          lut[11360] <= 16'd13580;
          lut[11361] <= 16'd13664;
          lut[11362] <= 16'd13748;
          lut[11363] <= 16'd13831;
          lut[11364] <= 16'd13912;
          lut[11365] <= 16'd13993;
          lut[11366] <= 16'd14073;
          lut[11367] <= 16'd14152;
          lut[11368] <= 16'd14230;
          lut[11369] <= 16'd14307;
          lut[11370] <= 16'd14384;
          lut[11371] <= 16'd14459;
          lut[11372] <= 16'd14534;
          lut[11373] <= 16'd14608;
          lut[11374] <= 16'd14681;
          lut[11375] <= 16'd14753;
          lut[11376] <= 16'd14825;
          lut[11377] <= 16'd14895;
          lut[11378] <= 16'd14965;
          lut[11379] <= 16'd15034;
          lut[11380] <= 16'd15103;
          lut[11381] <= 16'd15170;
          lut[11382] <= 16'd15237;
          lut[11383] <= 16'd15304;
          lut[11384] <= 16'd15369;
          lut[11385] <= 16'd15434;
          lut[11386] <= 16'd15498;
          lut[11387] <= 16'd15561;
          lut[11388] <= 16'd15624;
          lut[11389] <= 16'd15686;
          lut[11390] <= 16'd15747;
          lut[11391] <= 16'd15808;
          lut[11392] <= 0;
          lut[11393] <= 16'd184;
          lut[11394] <= 16'd368;
          lut[11395] <= 16'd552;
          lut[11396] <= 16'd736;
          lut[11397] <= 16'd919;
          lut[11398] <= 16'd1103;
          lut[11399] <= 16'd1286;
          lut[11400] <= 16'd1469;
          lut[11401] <= 16'd1651;
          lut[11402] <= 16'd1833;
          lut[11403] <= 16'd2015;
          lut[11404] <= 16'd2196;
          lut[11405] <= 16'd2376;
          lut[11406] <= 16'd2556;
          lut[11407] <= 16'd2736;
          lut[11408] <= 16'd2914;
          lut[11409] <= 16'd3092;
          lut[11410] <= 16'd3270;
          lut[11411] <= 16'd3446;
          lut[11412] <= 16'd3622;
          lut[11413] <= 16'd3796;
          lut[11414] <= 16'd3970;
          lut[11415] <= 16'd4143;
          lut[11416] <= 16'd4316;
          lut[11417] <= 16'd4487;
          lut[11418] <= 16'd4657;
          lut[11419] <= 16'd4826;
          lut[11420] <= 16'd4994;
          lut[11421] <= 16'd5161;
          lut[11422] <= 16'd5327;
          lut[11423] <= 16'd5491;
          lut[11424] <= 16'd5655;
          lut[11425] <= 16'd5817;
          lut[11426] <= 16'd5979;
          lut[11427] <= 16'd6139;
          lut[11428] <= 16'd6298;
          lut[11429] <= 16'd6455;
          lut[11430] <= 16'd6612;
          lut[11431] <= 16'd6767;
          lut[11432] <= 16'd6920;
          lut[11433] <= 16'd7073;
          lut[11434] <= 16'd7224;
          lut[11435] <= 16'd7374;
          lut[11436] <= 16'd7523;
          lut[11437] <= 16'd7670;
          lut[11438] <= 16'd7816;
          lut[11439] <= 16'd7960;
          lut[11440] <= 16'd8104;
          lut[11441] <= 16'd8246;
          lut[11442] <= 16'd8386;
          lut[11443] <= 16'd8526;
          lut[11444] <= 16'd8663;
          lut[11445] <= 16'd8800;
          lut[11446] <= 16'd8935;
          lut[11447] <= 16'd9069;
          lut[11448] <= 16'd9202;
          lut[11449] <= 16'd9333;
          lut[11450] <= 16'd9463;
          lut[11451] <= 16'd9591;
          lut[11452] <= 16'd9719;
          lut[11453] <= 16'd9844;
          lut[11454] <= 16'd9969;
          lut[11455] <= 16'd10092;
          lut[11456] <= 16'd10214;
          lut[11457] <= 16'd10335;
          lut[11458] <= 16'd10454;
          lut[11459] <= 16'd10573;
          lut[11460] <= 16'd10689;
          lut[11461] <= 16'd10805;
          lut[11462] <= 16'd10919;
          lut[11463] <= 16'd11032;
          lut[11464] <= 16'd11144;
          lut[11465] <= 16'd11255;
          lut[11466] <= 16'd11364;
          lut[11467] <= 16'd11473;
          lut[11468] <= 16'd11580;
          lut[11469] <= 16'd11686;
          lut[11470] <= 16'd11790;
          lut[11471] <= 16'd11894;
          lut[11472] <= 16'd11996;
          lut[11473] <= 16'd12098;
          lut[11474] <= 16'd12198;
          lut[11475] <= 16'd12297;
          lut[11476] <= 16'd12395;
          lut[11477] <= 16'd12491;
          lut[11478] <= 16'd12587;
          lut[11479] <= 16'd12682;
          lut[11480] <= 16'd12775;
          lut[11481] <= 16'd12868;
          lut[11482] <= 16'd12959;
          lut[11483] <= 16'd13050;
          lut[11484] <= 16'd13139;
          lut[11485] <= 16'd13228;
          lut[11486] <= 16'd13316;
          lut[11487] <= 16'd13402;
          lut[11488] <= 16'd13488;
          lut[11489] <= 16'd13572;
          lut[11490] <= 16'd13656;
          lut[11491] <= 16'd13739;
          lut[11492] <= 16'd13820;
          lut[11493] <= 16'd13901;
          lut[11494] <= 16'd13981;
          lut[11495] <= 16'd14061;
          lut[11496] <= 16'd14139;
          lut[11497] <= 16'd14216;
          lut[11498] <= 16'd14293;
          lut[11499] <= 16'd14368;
          lut[11500] <= 16'd14443;
          lut[11501] <= 16'd14517;
          lut[11502] <= 16'd14591;
          lut[11503] <= 16'd14663;
          lut[11504] <= 16'd14735;
          lut[11505] <= 16'd14805;
          lut[11506] <= 16'd14876;
          lut[11507] <= 16'd14945;
          lut[11508] <= 16'd15014;
          lut[11509] <= 16'd15081;
          lut[11510] <= 16'd15148;
          lut[11511] <= 16'd15215;
          lut[11512] <= 16'd15281;
          lut[11513] <= 16'd15346;
          lut[11514] <= 16'd15410;
          lut[11515] <= 16'd15473;
          lut[11516] <= 16'd15536;
          lut[11517] <= 16'd15599;
          lut[11518] <= 16'd15660;
          lut[11519] <= 16'd15721;
          lut[11520] <= 0;
          lut[11521] <= 16'd182;
          lut[11522] <= 16'd364;
          lut[11523] <= 16'd546;
          lut[11524] <= 16'd728;
          lut[11525] <= 16'd909;
          lut[11526] <= 16'd1091;
          lut[11527] <= 16'd1272;
          lut[11528] <= 16'd1453;
          lut[11529] <= 16'd1633;
          lut[11530] <= 16'd1813;
          lut[11531] <= 16'd1993;
          lut[11532] <= 16'd2172;
          lut[11533] <= 16'd2350;
          lut[11534] <= 16'd2528;
          lut[11535] <= 16'd2706;
          lut[11536] <= 16'd2883;
          lut[11537] <= 16'd3059;
          lut[11538] <= 16'd3234;
          lut[11539] <= 16'd3409;
          lut[11540] <= 16'd3583;
          lut[11541] <= 16'd3756;
          lut[11542] <= 16'd3928;
          lut[11543] <= 16'd4099;
          lut[11544] <= 16'd4270;
          lut[11545] <= 16'd4439;
          lut[11546] <= 16'd4608;
          lut[11547] <= 16'd4775;
          lut[11548] <= 16'd4942;
          lut[11549] <= 16'd5107;
          lut[11550] <= 16'd5272;
          lut[11551] <= 16'd5435;
          lut[11552] <= 16'd5597;
          lut[11553] <= 16'd5758;
          lut[11554] <= 16'd5918;
          lut[11555] <= 16'd6077;
          lut[11556] <= 16'd6234;
          lut[11557] <= 16'd6391;
          lut[11558] <= 16'd6546;
          lut[11559] <= 16'd6700;
          lut[11560] <= 16'd6852;
          lut[11561] <= 16'd7004;
          lut[11562] <= 16'd7154;
          lut[11563] <= 16'd7303;
          lut[11564] <= 16'd7450;
          lut[11565] <= 16'd7596;
          lut[11566] <= 16'd7741;
          lut[11567] <= 16'd7885;
          lut[11568] <= 16'd8027;
          lut[11569] <= 16'd8169;
          lut[11570] <= 16'd8308;
          lut[11571] <= 16'd8447;
          lut[11572] <= 16'd8584;
          lut[11573] <= 16'd8720;
          lut[11574] <= 16'd8854;
          lut[11575] <= 16'd8987;
          lut[11576] <= 16'd9119;
          lut[11577] <= 16'd9250;
          lut[11578] <= 16'd9379;
          lut[11579] <= 16'd9507;
          lut[11580] <= 16'd9634;
          lut[11581] <= 16'd9759;
          lut[11582] <= 16'd9883;
          lut[11583] <= 16'd10006;
          lut[11584] <= 16'd10128;
          lut[11585] <= 16'd10248;
          lut[11586] <= 16'd10367;
          lut[11587] <= 16'd10485;
          lut[11588] <= 16'd10601;
          lut[11589] <= 16'd10716;
          lut[11590] <= 16'd10831;
          lut[11591] <= 16'd10943;
          lut[11592] <= 16'd11055;
          lut[11593] <= 16'd11165;
          lut[11594] <= 16'd11275;
          lut[11595] <= 16'd11383;
          lut[11596] <= 16'd11489;
          lut[11597] <= 16'd11595;
          lut[11598] <= 16'd11700;
          lut[11599] <= 16'd11803;
          lut[11600] <= 16'd11905;
          lut[11601] <= 16'd12006;
          lut[11602] <= 16'd12106;
          lut[11603] <= 16'd12205;
          lut[11604] <= 16'd12303;
          lut[11605] <= 16'd12400;
          lut[11606] <= 16'd12496;
          lut[11607] <= 16'd12590;
          lut[11608] <= 16'd12684;
          lut[11609] <= 16'd12776;
          lut[11610] <= 16'd12868;
          lut[11611] <= 16'd12958;
          lut[11612] <= 16'd13048;
          lut[11613] <= 16'd13137;
          lut[11614] <= 16'd13224;
          lut[11615] <= 16'd13311;
          lut[11616] <= 16'd13396;
          lut[11617] <= 16'd13481;
          lut[11618] <= 16'd13565;
          lut[11619] <= 16'd13648;
          lut[11620] <= 16'd13729;
          lut[11621] <= 16'd13811;
          lut[11622] <= 16'd13891;
          lut[11623] <= 16'd13970;
          lut[11624] <= 16'd14048;
          lut[11625] <= 16'd14126;
          lut[11626] <= 16'd14202;
          lut[11627] <= 16'd14278;
          lut[11628] <= 16'd14353;
          lut[11629] <= 16'd14428;
          lut[11630] <= 16'd14501;
          lut[11631] <= 16'd14574;
          lut[11632] <= 16'd14645;
          lut[11633] <= 16'd14716;
          lut[11634] <= 16'd14787;
          lut[11635] <= 16'd14856;
          lut[11636] <= 16'd14925;
          lut[11637] <= 16'd14993;
          lut[11638] <= 16'd15060;
          lut[11639] <= 16'd15127;
          lut[11640] <= 16'd15193;
          lut[11641] <= 16'd15258;
          lut[11642] <= 16'd15322;
          lut[11643] <= 16'd15386;
          lut[11644] <= 16'd15449;
          lut[11645] <= 16'd15512;
          lut[11646] <= 16'd15574;
          lut[11647] <= 16'd15635;
          lut[11648] <= 0;
          lut[11649] <= 16'd180;
          lut[11650] <= 16'd360;
          lut[11651] <= 16'd540;
          lut[11652] <= 16'd720;
          lut[11653] <= 16'd899;
          lut[11654] <= 16'd1079;
          lut[11655] <= 16'd1258;
          lut[11656] <= 16'd1437;
          lut[11657] <= 16'd1615;
          lut[11658] <= 16'd1793;
          lut[11659] <= 16'd1971;
          lut[11660] <= 16'd2148;
          lut[11661] <= 16'd2325;
          lut[11662] <= 16'd2501;
          lut[11663] <= 16'd2677;
          lut[11664] <= 16'd2852;
          lut[11665] <= 16'd3026;
          lut[11666] <= 16'd3199;
          lut[11667] <= 16'd3372;
          lut[11668] <= 16'd3545;
          lut[11669] <= 16'd3716;
          lut[11670] <= 16'd3886;
          lut[11671] <= 16'd4056;
          lut[11672] <= 16'd4225;
          lut[11673] <= 16'd4393;
          lut[11674] <= 16'd4560;
          lut[11675] <= 16'd4726;
          lut[11676] <= 16'd4891;
          lut[11677] <= 16'd5055;
          lut[11678] <= 16'd5217;
          lut[11679] <= 16'd5379;
          lut[11680] <= 16'd5540;
          lut[11681] <= 16'd5700;
          lut[11682] <= 16'd5858;
          lut[11683] <= 16'd6016;
          lut[11684] <= 16'd6172;
          lut[11685] <= 16'd6327;
          lut[11686] <= 16'd6481;
          lut[11687] <= 16'd6634;
          lut[11688] <= 16'd6785;
          lut[11689] <= 16'd6936;
          lut[11690] <= 16'd7085;
          lut[11691] <= 16'd7232;
          lut[11692] <= 16'd7379;
          lut[11693] <= 16'd7524;
          lut[11694] <= 16'd7668;
          lut[11695] <= 16'd7811;
          lut[11696] <= 16'd7953;
          lut[11697] <= 16'd8093;
          lut[11698] <= 16'd8232;
          lut[11699] <= 16'd8369;
          lut[11700] <= 16'd8506;
          lut[11701] <= 16'd8641;
          lut[11702] <= 16'd8775;
          lut[11703] <= 16'd8907;
          lut[11704] <= 16'd9038;
          lut[11705] <= 16'd9168;
          lut[11706] <= 16'd9297;
          lut[11707] <= 16'd9424;
          lut[11708] <= 16'd9550;
          lut[11709] <= 16'd9675;
          lut[11710] <= 16'd9799;
          lut[11711] <= 16'd9921;
          lut[11712] <= 16'd10042;
          lut[11713] <= 16'd10162;
          lut[11714] <= 16'd10281;
          lut[11715] <= 16'd10398;
          lut[11716] <= 16'd10514;
          lut[11717] <= 16'd10629;
          lut[11718] <= 16'd10743;
          lut[11719] <= 16'd10855;
          lut[11720] <= 16'd10967;
          lut[11721] <= 16'd11077;
          lut[11722] <= 16'd11186;
          lut[11723] <= 16'd11294;
          lut[11724] <= 16'd11400;
          lut[11725] <= 16'd11506;
          lut[11726] <= 16'd11610;
          lut[11727] <= 16'd11713;
          lut[11728] <= 16'd11815;
          lut[11729] <= 16'd11916;
          lut[11730] <= 16'd12016;
          lut[11731] <= 16'd12115;
          lut[11732] <= 16'd12213;
          lut[11733] <= 16'd12310;
          lut[11734] <= 16'd12405;
          lut[11735] <= 16'd12500;
          lut[11736] <= 16'd12593;
          lut[11737] <= 16'd12686;
          lut[11738] <= 16'd12777;
          lut[11739] <= 16'd12868;
          lut[11740] <= 16'd12957;
          lut[11741] <= 16'd13046;
          lut[11742] <= 16'd13134;
          lut[11743] <= 16'd13220;
          lut[11744] <= 16'd13306;
          lut[11745] <= 16'd13391;
          lut[11746] <= 16'd13475;
          lut[11747] <= 16'd13557;
          lut[11748] <= 16'd13639;
          lut[11749] <= 16'd13721;
          lut[11750] <= 16'd13801;
          lut[11751] <= 16'd13880;
          lut[11752] <= 16'd13959;
          lut[11753] <= 16'd14036;
          lut[11754] <= 16'd14113;
          lut[11755] <= 16'd14189;
          lut[11756] <= 16'd14264;
          lut[11757] <= 16'd14339;
          lut[11758] <= 16'd14412;
          lut[11759] <= 16'd14485;
          lut[11760] <= 16'd14557;
          lut[11761] <= 16'd14628;
          lut[11762] <= 16'd14699;
          lut[11763] <= 16'd14768;
          lut[11764] <= 16'd14837;
          lut[11765] <= 16'd14905;
          lut[11766] <= 16'd14973;
          lut[11767] <= 16'd15040;
          lut[11768] <= 16'd15106;
          lut[11769] <= 16'd15171;
          lut[11770] <= 16'd15236;
          lut[11771] <= 16'd15300;
          lut[11772] <= 16'd15363;
          lut[11773] <= 16'd15426;
          lut[11774] <= 16'd15488;
          lut[11775] <= 16'd15549;
          lut[11776] <= 0;
          lut[11777] <= 16'd178;
          lut[11778] <= 16'd356;
          lut[11779] <= 16'd534;
          lut[11780] <= 16'd712;
          lut[11781] <= 16'd890;
          lut[11782] <= 16'd1067;
          lut[11783] <= 16'd1244;
          lut[11784] <= 16'd1421;
          lut[11785] <= 16'd1598;
          lut[11786] <= 16'd1774;
          lut[11787] <= 16'd1950;
          lut[11788] <= 16'd2125;
          lut[11789] <= 16'd2300;
          lut[11790] <= 16'd2474;
          lut[11791] <= 16'd2648;
          lut[11792] <= 16'd2821;
          lut[11793] <= 16'd2994;
          lut[11794] <= 16'd3166;
          lut[11795] <= 16'd3337;
          lut[11796] <= 16'd3507;
          lut[11797] <= 16'd3677;
          lut[11798] <= 16'd3846;
          lut[11799] <= 16'd4014;
          lut[11800] <= 16'd4181;
          lut[11801] <= 16'd4347;
          lut[11802] <= 16'd4513;
          lut[11803] <= 16'd4677;
          lut[11804] <= 16'd4841;
          lut[11805] <= 16'd5003;
          lut[11806] <= 16'd5164;
          lut[11807] <= 16'd5325;
          lut[11808] <= 16'd5484;
          lut[11809] <= 16'd5643;
          lut[11810] <= 16'd5800;
          lut[11811] <= 16'd5956;
          lut[11812] <= 16'd6111;
          lut[11813] <= 16'd6265;
          lut[11814] <= 16'd6418;
          lut[11815] <= 16'd6569;
          lut[11816] <= 16'd6720;
          lut[11817] <= 16'd6869;
          lut[11818] <= 16'd7017;
          lut[11819] <= 16'd7163;
          lut[11820] <= 16'd7309;
          lut[11821] <= 16'd7453;
          lut[11822] <= 16'd7596;
          lut[11823] <= 16'd7738;
          lut[11824] <= 16'd7879;
          lut[11825] <= 16'd8018;
          lut[11826] <= 16'd8156;
          lut[11827] <= 16'd8293;
          lut[11828] <= 16'd8429;
          lut[11829] <= 16'd8563;
          lut[11830] <= 16'd8696;
          lut[11831] <= 16'd8828;
          lut[11832] <= 16'd8959;
          lut[11833] <= 16'd9088;
          lut[11834] <= 16'd9216;
          lut[11835] <= 16'd9343;
          lut[11836] <= 16'd9468;
          lut[11837] <= 16'd9593;
          lut[11838] <= 16'd9716;
          lut[11839] <= 16'd9838;
          lut[11840] <= 16'd9958;
          lut[11841] <= 16'd10078;
          lut[11842] <= 16'd10196;
          lut[11843] <= 16'd10313;
          lut[11844] <= 16'd10429;
          lut[11845] <= 16'd10543;
          lut[11846] <= 16'd10657;
          lut[11847] <= 16'd10769;
          lut[11848] <= 16'd10880;
          lut[11849] <= 16'd10990;
          lut[11850] <= 16'd11098;
          lut[11851] <= 16'd11206;
          lut[11852] <= 16'd11312;
          lut[11853] <= 16'd11418;
          lut[11854] <= 16'd11522;
          lut[11855] <= 16'd11625;
          lut[11856] <= 16'd11727;
          lut[11857] <= 16'd11828;
          lut[11858] <= 16'd11927;
          lut[11859] <= 16'd12026;
          lut[11860] <= 16'd12124;
          lut[11861] <= 16'd12220;
          lut[11862] <= 16'd12316;
          lut[11863] <= 16'd12410;
          lut[11864] <= 16'd12504;
          lut[11865] <= 16'd12596;
          lut[11866] <= 16'd12688;
          lut[11867] <= 16'd12778;
          lut[11868] <= 16'd12868;
          lut[11869] <= 16'd12957;
          lut[11870] <= 16'd13044;
          lut[11871] <= 16'd13131;
          lut[11872] <= 16'd13217;
          lut[11873] <= 16'd13301;
          lut[11874] <= 16'd13385;
          lut[11875] <= 16'd13468;
          lut[11876] <= 16'd13550;
          lut[11877] <= 16'd13631;
          lut[11878] <= 16'd13712;
          lut[11879] <= 16'd13791;
          lut[11880] <= 16'd13870;
          lut[11881] <= 16'd13948;
          lut[11882] <= 16'd14025;
          lut[11883] <= 16'd14101;
          lut[11884] <= 16'd14176;
          lut[11885] <= 16'd14250;
          lut[11886] <= 16'd14324;
          lut[11887] <= 16'd14397;
          lut[11888] <= 16'd14469;
          lut[11889] <= 16'd14540;
          lut[11890] <= 16'd14611;
          lut[11891] <= 16'd14681;
          lut[11892] <= 16'd14750;
          lut[11893] <= 16'd14819;
          lut[11894] <= 16'd14886;
          lut[11895] <= 16'd14953;
          lut[11896] <= 16'd15019;
          lut[11897] <= 16'd15085;
          lut[11898] <= 16'd15150;
          lut[11899] <= 16'd15214;
          lut[11900] <= 16'd15278;
          lut[11901] <= 16'd15341;
          lut[11902] <= 16'd15403;
          lut[11903] <= 16'd15464;
          lut[11904] <= 0;
          lut[11905] <= 16'd176;
          lut[11906] <= 16'd352;
          lut[11907] <= 16'd528;
          lut[11908] <= 16'd704;
          lut[11909] <= 16'd880;
          lut[11910] <= 16'd1056;
          lut[11911] <= 16'd1231;
          lut[11912] <= 16'd1406;
          lut[11913] <= 16'd1581;
          lut[11914] <= 16'd1755;
          lut[11915] <= 16'd1929;
          lut[11916] <= 16'd2102;
          lut[11917] <= 16'd2275;
          lut[11918] <= 16'd2448;
          lut[11919] <= 16'd2620;
          lut[11920] <= 16'd2791;
          lut[11921] <= 16'd2962;
          lut[11922] <= 16'd3132;
          lut[11923] <= 16'd3302;
          lut[11924] <= 16'd3471;
          lut[11925] <= 16'd3639;
          lut[11926] <= 16'd3806;
          lut[11927] <= 16'd3972;
          lut[11928] <= 16'd4138;
          lut[11929] <= 16'd4303;
          lut[11930] <= 16'd4466;
          lut[11931] <= 16'd4629;
          lut[11932] <= 16'd4791;
          lut[11933] <= 16'd4952;
          lut[11934] <= 16'd5112;
          lut[11935] <= 16'd5272;
          lut[11936] <= 16'd5430;
          lut[11937] <= 16'd5587;
          lut[11938] <= 16'd5743;
          lut[11939] <= 16'd5897;
          lut[11940] <= 16'd6051;
          lut[11941] <= 16'd6204;
          lut[11942] <= 16'd6355;
          lut[11943] <= 16'd6506;
          lut[11944] <= 16'd6655;
          lut[11945] <= 16'd6803;
          lut[11946] <= 16'd6950;
          lut[11947] <= 16'd7096;
          lut[11948] <= 16'd7240;
          lut[11949] <= 16'd7384;
          lut[11950] <= 16'd7526;
          lut[11951] <= 16'd7667;
          lut[11952] <= 16'd7806;
          lut[11953] <= 16'd7945;
          lut[11954] <= 16'd8082;
          lut[11955] <= 16'd8218;
          lut[11956] <= 16'd8353;
          lut[11957] <= 16'd8487;
          lut[11958] <= 16'd8619;
          lut[11959] <= 16'd8750;
          lut[11960] <= 16'd8880;
          lut[11961] <= 16'd9009;
          lut[11962] <= 16'd9136;
          lut[11963] <= 16'd9262;
          lut[11964] <= 16'd9387;
          lut[11965] <= 16'd9511;
          lut[11966] <= 16'd9634;
          lut[11967] <= 16'd9755;
          lut[11968] <= 16'd9875;
          lut[11969] <= 16'd9994;
          lut[11970] <= 16'd10112;
          lut[11971] <= 16'd10229;
          lut[11972] <= 16'd10344;
          lut[11973] <= 16'd10458;
          lut[11974] <= 16'd10571;
          lut[11975] <= 16'd10683;
          lut[11976] <= 16'd10794;
          lut[11977] <= 16'd10903;
          lut[11978] <= 16'd11012;
          lut[11979] <= 16'd11119;
          lut[11980] <= 16'd11225;
          lut[11981] <= 16'd11330;
          lut[11982] <= 16'd11434;
          lut[11983] <= 16'd11537;
          lut[11984] <= 16'd11639;
          lut[11985] <= 16'd11740;
          lut[11986] <= 16'd11839;
          lut[11987] <= 16'd11938;
          lut[11988] <= 16'd12036;
          lut[11989] <= 16'd12132;
          lut[11990] <= 16'd12228;
          lut[11991] <= 16'd12322;
          lut[11992] <= 16'd12415;
          lut[11993] <= 16'd12508;
          lut[11994] <= 16'd12599;
          lut[11995] <= 16'd12690;
          lut[11996] <= 16'd12779;
          lut[11997] <= 16'd12868;
          lut[11998] <= 16'd12956;
          lut[11999] <= 16'd13042;
          lut[12000] <= 16'd13128;
          lut[12001] <= 16'd13213;
          lut[12002] <= 16'd13297;
          lut[12003] <= 16'd13380;
          lut[12004] <= 16'd13462;
          lut[12005] <= 16'd13543;
          lut[12006] <= 16'd13624;
          lut[12007] <= 16'd13703;
          lut[12008] <= 16'd13782;
          lut[12009] <= 16'd13860;
          lut[12010] <= 16'd13937;
          lut[12011] <= 16'd14013;
          lut[12012] <= 16'd14088;
          lut[12013] <= 16'd14163;
          lut[12014] <= 16'd14237;
          lut[12015] <= 16'd14310;
          lut[12016] <= 16'd14382;
          lut[12017] <= 16'd14454;
          lut[12018] <= 16'd14524;
          lut[12019] <= 16'd14594;
          lut[12020] <= 16'd14664;
          lut[12021] <= 16'd14732;
          lut[12022] <= 16'd14800;
          lut[12023] <= 16'd14867;
          lut[12024] <= 16'd14934;
          lut[12025] <= 16'd15000;
          lut[12026] <= 16'd15065;
          lut[12027] <= 16'd15129;
          lut[12028] <= 16'd15193;
          lut[12029] <= 16'd15256;
          lut[12030] <= 16'd15318;
          lut[12031] <= 16'd15380;
          lut[12032] <= 0;
          lut[12033] <= 16'd174;
          lut[12034] <= 16'd349;
          lut[12035] <= 16'd523;
          lut[12036] <= 16'd697;
          lut[12037] <= 16'd871;
          lut[12038] <= 16'd1044;
          lut[12039] <= 16'd1218;
          lut[12040] <= 16'd1391;
          lut[12041] <= 16'd1564;
          lut[12042] <= 16'd1736;
          lut[12043] <= 16'd1909;
          lut[12044] <= 16'd2080;
          lut[12045] <= 16'd2252;
          lut[12046] <= 16'd2422;
          lut[12047] <= 16'd2593;
          lut[12048] <= 16'd2762;
          lut[12049] <= 16'd2931;
          lut[12050] <= 16'd3100;
          lut[12051] <= 16'd3268;
          lut[12052] <= 16'd3435;
          lut[12053] <= 16'd3601;
          lut[12054] <= 16'd3767;
          lut[12055] <= 16'd3932;
          lut[12056] <= 16'd4096;
          lut[12057] <= 16'd4259;
          lut[12058] <= 16'd4421;
          lut[12059] <= 16'd4583;
          lut[12060] <= 16'd4743;
          lut[12061] <= 16'd4903;
          lut[12062] <= 16'd5062;
          lut[12063] <= 16'd5219;
          lut[12064] <= 16'd5376;
          lut[12065] <= 16'd5532;
          lut[12066] <= 16'd5686;
          lut[12067] <= 16'd5840;
          lut[12068] <= 16'd5992;
          lut[12069] <= 16'd6144;
          lut[12070] <= 16'd6294;
          lut[12071] <= 16'd6443;
          lut[12072] <= 16'd6592;
          lut[12073] <= 16'd6739;
          lut[12074] <= 16'd6885;
          lut[12075] <= 16'd7029;
          lut[12076] <= 16'd7173;
          lut[12077] <= 16'd7315;
          lut[12078] <= 16'd7456;
          lut[12079] <= 16'd7596;
          lut[12080] <= 16'd7735;
          lut[12081] <= 16'd7873;
          lut[12082] <= 16'd8009;
          lut[12083] <= 16'd8145;
          lut[12084] <= 16'd8279;
          lut[12085] <= 16'd8412;
          lut[12086] <= 16'd8543;
          lut[12087] <= 16'd8674;
          lut[12088] <= 16'd8803;
          lut[12089] <= 16'd8931;
          lut[12090] <= 16'd9058;
          lut[12091] <= 16'd9183;
          lut[12092] <= 16'd9308;
          lut[12093] <= 16'd9431;
          lut[12094] <= 16'd9553;
          lut[12095] <= 16'd9674;
          lut[12096] <= 16'd9794;
          lut[12097] <= 16'd9912;
          lut[12098] <= 16'd10030;
          lut[12099] <= 16'd10146;
          lut[12100] <= 16'd10261;
          lut[12101] <= 16'd10375;
          lut[12102] <= 16'd10487;
          lut[12103] <= 16'd10599;
          lut[12104] <= 16'd10709;
          lut[12105] <= 16'd10818;
          lut[12106] <= 16'd10927;
          lut[12107] <= 16'd11034;
          lut[12108] <= 16'd11140;
          lut[12109] <= 16'd11244;
          lut[12110] <= 16'd11348;
          lut[12111] <= 16'd11451;
          lut[12112] <= 16'd11553;
          lut[12113] <= 16'd11653;
          lut[12114] <= 16'd11753;
          lut[12115] <= 16'd11851;
          lut[12116] <= 16'd11948;
          lut[12117] <= 16'd12045;
          lut[12118] <= 16'd12140;
          lut[12119] <= 16'd12235;
          lut[12120] <= 16'd12328;
          lut[12121] <= 16'd12420;
          lut[12122] <= 16'd12512;
          lut[12123] <= 16'd12602;
          lut[12124] <= 16'd12692;
          lut[12125] <= 16'd12780;
          lut[12126] <= 16'd12868;
          lut[12127] <= 16'd12955;
          lut[12128] <= 16'd13040;
          lut[12129] <= 16'd13125;
          lut[12130] <= 16'd13209;
          lut[12131] <= 16'd13292;
          lut[12132] <= 16'd13375;
          lut[12133] <= 16'd13456;
          lut[12134] <= 16'd13536;
          lut[12135] <= 16'd13616;
          lut[12136] <= 16'd13695;
          lut[12137] <= 16'd13773;
          lut[12138] <= 16'd13850;
          lut[12139] <= 16'd13926;
          lut[12140] <= 16'd14002;
          lut[12141] <= 16'd14076;
          lut[12142] <= 16'd14150;
          lut[12143] <= 16'd14224;
          lut[12144] <= 16'd14296;
          lut[12145] <= 16'd14368;
          lut[12146] <= 16'd14439;
          lut[12147] <= 16'd14509;
          lut[12148] <= 16'd14578;
          lut[12149] <= 16'd14647;
          lut[12150] <= 16'd14715;
          lut[12151] <= 16'd14782;
          lut[12152] <= 16'd14849;
          lut[12153] <= 16'd14915;
          lut[12154] <= 16'd14980;
          lut[12155] <= 16'd15045;
          lut[12156] <= 16'd15109;
          lut[12157] <= 16'd15172;
          lut[12158] <= 16'd15234;
          lut[12159] <= 16'd15296;
          lut[12160] <= 0;
          lut[12161] <= 16'd172;
          lut[12162] <= 16'd345;
          lut[12163] <= 16'd517;
          lut[12164] <= 16'd689;
          lut[12165] <= 16'd862;
          lut[12166] <= 16'd1033;
          lut[12167] <= 16'd1205;
          lut[12168] <= 16'd1376;
          lut[12169] <= 16'd1548;
          lut[12170] <= 16'd1718;
          lut[12171] <= 16'd1889;
          lut[12172] <= 16'd2059;
          lut[12173] <= 16'd2228;
          lut[12174] <= 16'd2397;
          lut[12175] <= 16'd2566;
          lut[12176] <= 16'd2734;
          lut[12177] <= 16'd2901;
          lut[12178] <= 16'd3068;
          lut[12179] <= 16'd3234;
          lut[12180] <= 16'd3400;
          lut[12181] <= 16'd3564;
          lut[12182] <= 16'd3728;
          lut[12183] <= 16'd3892;
          lut[12184] <= 16'd4054;
          lut[12185] <= 16'd4216;
          lut[12186] <= 16'd4377;
          lut[12187] <= 16'd4537;
          lut[12188] <= 16'd4696;
          lut[12189] <= 16'd4854;
          lut[12190] <= 16'd5012;
          lut[12191] <= 16'd5168;
          lut[12192] <= 16'd5323;
          lut[12193] <= 16'd5478;
          lut[12194] <= 16'd5631;
          lut[12195] <= 16'd5783;
          lut[12196] <= 16'd5935;
          lut[12197] <= 16'd6085;
          lut[12198] <= 16'd6234;
          lut[12199] <= 16'd6382;
          lut[12200] <= 16'd6529;
          lut[12201] <= 16'd6675;
          lut[12202] <= 16'd6820;
          lut[12203] <= 16'd6964;
          lut[12204] <= 16'd7106;
          lut[12205] <= 16'd7248;
          lut[12206] <= 16'd7388;
          lut[12207] <= 16'd7527;
          lut[12208] <= 16'd7665;
          lut[12209] <= 16'd7802;
          lut[12210] <= 16'd7938;
          lut[12211] <= 16'd8072;
          lut[12212] <= 16'd8205;
          lut[12213] <= 16'd8338;
          lut[12214] <= 16'd8468;
          lut[12215] <= 16'd8598;
          lut[12216] <= 16'd8727;
          lut[12217] <= 16'd8854;
          lut[12218] <= 16'd8980;
          lut[12219] <= 16'd9106;
          lut[12220] <= 16'd9229;
          lut[12221] <= 16'd9352;
          lut[12222] <= 16'd9474;
          lut[12223] <= 16'd9594;
          lut[12224] <= 16'd9713;
          lut[12225] <= 16'd9831;
          lut[12226] <= 16'd9948;
          lut[12227] <= 16'd10064;
          lut[12228] <= 16'd10178;
          lut[12229] <= 16'd10292;
          lut[12230] <= 16'd10404;
          lut[12231] <= 16'd10515;
          lut[12232] <= 16'd10626;
          lut[12233] <= 16'd10735;
          lut[12234] <= 16'd10842;
          lut[12235] <= 16'd10949;
          lut[12236] <= 16'd11055;
          lut[12237] <= 16'd11160;
          lut[12238] <= 16'd11263;
          lut[12239] <= 16'd11366;
          lut[12240] <= 16'd11467;
          lut[12241] <= 16'd11567;
          lut[12242] <= 16'd11667;
          lut[12243] <= 16'd11765;
          lut[12244] <= 16'd11862;
          lut[12245] <= 16'd11959;
          lut[12246] <= 16'd12054;
          lut[12247] <= 16'd12148;
          lut[12248] <= 16'd12242;
          lut[12249] <= 16'd12334;
          lut[12250] <= 16'd12425;
          lut[12251] <= 16'd12516;
          lut[12252] <= 16'd12605;
          lut[12253] <= 16'd12694;
          lut[12254] <= 16'd12781;
          lut[12255] <= 16'd12868;
          lut[12256] <= 16'd12954;
          lut[12257] <= 16'd13039;
          lut[12258] <= 16'd13123;
          lut[12259] <= 16'd13206;
          lut[12260] <= 16'd13288;
          lut[12261] <= 16'd13369;
          lut[12262] <= 16'd13450;
          lut[12263] <= 16'd13530;
          lut[12264] <= 16'd13608;
          lut[12265] <= 16'd13686;
          lut[12266] <= 16'd13764;
          lut[12267] <= 16'd13840;
          lut[12268] <= 16'd13916;
          lut[12269] <= 16'd13991;
          lut[12270] <= 16'd14065;
          lut[12271] <= 16'd14138;
          lut[12272] <= 16'd14210;
          lut[12273] <= 16'd14282;
          lut[12274] <= 16'd14353;
          lut[12275] <= 16'd14424;
          lut[12276] <= 16'd14493;
          lut[12277] <= 16'd14562;
          lut[12278] <= 16'd14630;
          lut[12279] <= 16'd14698;
          lut[12280] <= 16'd14765;
          lut[12281] <= 16'd14831;
          lut[12282] <= 16'd14896;
          lut[12283] <= 16'd14961;
          lut[12284] <= 16'd15025;
          lut[12285] <= 16'd15088;
          lut[12286] <= 16'd15151;
          lut[12287] <= 16'd15213;
          lut[12288] <= 0;
          lut[12289] <= 16'd171;
          lut[12290] <= 16'd341;
          lut[12291] <= 16'd512;
          lut[12292] <= 16'd682;
          lut[12293] <= 16'd853;
          lut[12294] <= 16'd1023;
          lut[12295] <= 16'd1193;
          lut[12296] <= 16'd1362;
          lut[12297] <= 16'd1532;
          lut[12298] <= 16'd1701;
          lut[12299] <= 16'd1869;
          lut[12300] <= 16'd2037;
          lut[12301] <= 16'd2205;
          lut[12302] <= 16'd2373;
          lut[12303] <= 16'd2539;
          lut[12304] <= 16'd2706;
          lut[12305] <= 16'd2872;
          lut[12306] <= 16'd3037;
          lut[12307] <= 16'd3201;
          lut[12308] <= 16'd3365;
          lut[12309] <= 16'd3528;
          lut[12310] <= 16'd3691;
          lut[12311] <= 16'd3853;
          lut[12312] <= 16'd4014;
          lut[12313] <= 16'd4174;
          lut[12314] <= 16'd4333;
          lut[12315] <= 16'd4492;
          lut[12316] <= 16'd4650;
          lut[12317] <= 16'd4807;
          lut[12318] <= 16'd4962;
          lut[12319] <= 16'd5117;
          lut[12320] <= 16'd5272;
          lut[12321] <= 16'd5425;
          lut[12322] <= 16'd5577;
          lut[12323] <= 16'd5728;
          lut[12324] <= 16'd5878;
          lut[12325] <= 16'd6027;
          lut[12326] <= 16'd6175;
          lut[12327] <= 16'd6322;
          lut[12328] <= 16'd6468;
          lut[12329] <= 16'd6613;
          lut[12330] <= 16'd6757;
          lut[12331] <= 16'd6900;
          lut[12332] <= 16'd7041;
          lut[12333] <= 16'd7182;
          lut[12334] <= 16'd7321;
          lut[12335] <= 16'd7459;
          lut[12336] <= 16'd7596;
          lut[12337] <= 16'd7732;
          lut[12338] <= 16'd7867;
          lut[12339] <= 16'd8001;
          lut[12340] <= 16'd8133;
          lut[12341] <= 16'd8265;
          lut[12342] <= 16'd8395;
          lut[12343] <= 16'd8524;
          lut[12344] <= 16'd8652;
          lut[12345] <= 16'd8779;
          lut[12346] <= 16'd8904;
          lut[12347] <= 16'd9029;
          lut[12348] <= 16'd9152;
          lut[12349] <= 16'd9274;
          lut[12350] <= 16'd9395;
          lut[12351] <= 16'd9515;
          lut[12352] <= 16'd9634;
          lut[12353] <= 16'd9751;
          lut[12354] <= 16'd9868;
          lut[12355] <= 16'd9983;
          lut[12356] <= 16'd10097;
          lut[12357] <= 16'd10210;
          lut[12358] <= 16'd10322;
          lut[12359] <= 16'd10433;
          lut[12360] <= 16'd10543;
          lut[12361] <= 16'd10652;
          lut[12362] <= 16'd10759;
          lut[12363] <= 16'd10866;
          lut[12364] <= 16'd10971;
          lut[12365] <= 16'd11076;
          lut[12366] <= 16'd11179;
          lut[12367] <= 16'd11281;
          lut[12368] <= 16'd11383;
          lut[12369] <= 16'd11483;
          lut[12370] <= 16'd11582;
          lut[12371] <= 16'd11680;
          lut[12372] <= 16'd11777;
          lut[12373] <= 16'd11873;
          lut[12374] <= 16'd11969;
          lut[12375] <= 16'd12063;
          lut[12376] <= 16'd12156;
          lut[12377] <= 16'd12248;
          lut[12378] <= 16'd12340;
          lut[12379] <= 16'd12430;
          lut[12380] <= 16'd12519;
          lut[12381] <= 16'd12608;
          lut[12382] <= 16'd12696;
          lut[12383] <= 16'd12782;
          lut[12384] <= 16'd12868;
          lut[12385] <= 16'd12953;
          lut[12386] <= 16'd13037;
          lut[12387] <= 16'd13120;
          lut[12388] <= 16'd13202;
          lut[12389] <= 16'd13284;
          lut[12390] <= 16'd13364;
          lut[12391] <= 16'd13444;
          lut[12392] <= 16'd13523;
          lut[12393] <= 16'd13601;
          lut[12394] <= 16'd13678;
          lut[12395] <= 16'd13755;
          lut[12396] <= 16'd13831;
          lut[12397] <= 16'd13906;
          lut[12398] <= 16'd13980;
          lut[12399] <= 16'd14053;
          lut[12400] <= 16'd14126;
          lut[12401] <= 16'd14198;
          lut[12402] <= 16'd14269;
          lut[12403] <= 16'd14339;
          lut[12404] <= 16'd14409;
          lut[12405] <= 16'd14478;
          lut[12406] <= 16'd14546;
          lut[12407] <= 16'd14614;
          lut[12408] <= 16'd14681;
          lut[12409] <= 16'd14747;
          lut[12410] <= 16'd14813;
          lut[12411] <= 16'd14878;
          lut[12412] <= 16'd14942;
          lut[12413] <= 16'd15006;
          lut[12414] <= 16'd15069;
          lut[12415] <= 16'd15131;
          lut[12416] <= 0;
          lut[12417] <= 16'd169;
          lut[12418] <= 16'd338;
          lut[12419] <= 16'd507;
          lut[12420] <= 16'd675;
          lut[12421] <= 16'd844;
          lut[12422] <= 16'd1012;
          lut[12423] <= 16'd1180;
          lut[12424] <= 16'd1348;
          lut[12425] <= 16'd1516;
          lut[12426] <= 16'd1683;
          lut[12427] <= 16'd1850;
          lut[12428] <= 16'd2017;
          lut[12429] <= 16'd2183;
          lut[12430] <= 16'd2348;
          lut[12431] <= 16'd2514;
          lut[12432] <= 16'd2678;
          lut[12433] <= 16'd2843;
          lut[12434] <= 16'd3006;
          lut[12435] <= 16'd3169;
          lut[12436] <= 16'd3331;
          lut[12437] <= 16'd3493;
          lut[12438] <= 16'd3654;
          lut[12439] <= 16'd3814;
          lut[12440] <= 16'd3974;
          lut[12441] <= 16'd4133;
          lut[12442] <= 16'd4291;
          lut[12443] <= 16'd4448;
          lut[12444] <= 16'd4604;
          lut[12445] <= 16'd4760;
          lut[12446] <= 16'd4914;
          lut[12447] <= 16'd5068;
          lut[12448] <= 16'd5221;
          lut[12449] <= 16'd5373;
          lut[12450] <= 16'd5524;
          lut[12451] <= 16'd5674;
          lut[12452] <= 16'd5822;
          lut[12453] <= 16'd5970;
          lut[12454] <= 16'd6117;
          lut[12455] <= 16'd6263;
          lut[12456] <= 16'd6408;
          lut[12457] <= 16'd6552;
          lut[12458] <= 16'd6695;
          lut[12459] <= 16'd6837;
          lut[12460] <= 16'd6977;
          lut[12461] <= 16'd7117;
          lut[12462] <= 16'd7255;
          lut[12463] <= 16'd7392;
          lut[12464] <= 16'd7529;
          lut[12465] <= 16'd7664;
          lut[12466] <= 16'd7798;
          lut[12467] <= 16'd7931;
          lut[12468] <= 16'd8062;
          lut[12469] <= 16'd8193;
          lut[12470] <= 16'd8323;
          lut[12471] <= 16'd8451;
          lut[12472] <= 16'd8578;
          lut[12473] <= 16'd8704;
          lut[12474] <= 16'd8829;
          lut[12475] <= 16'd8953;
          lut[12476] <= 16'd9076;
          lut[12477] <= 16'd9198;
          lut[12478] <= 16'd9318;
          lut[12479] <= 16'd9437;
          lut[12480] <= 16'd9556;
          lut[12481] <= 16'd9673;
          lut[12482] <= 16'd9789;
          lut[12483] <= 16'd9904;
          lut[12484] <= 16'd10017;
          lut[12485] <= 16'd10130;
          lut[12486] <= 16'd10242;
          lut[12487] <= 16'd10352;
          lut[12488] <= 16'd10462;
          lut[12489] <= 16'd10570;
          lut[12490] <= 16'd10677;
          lut[12491] <= 16'd10784;
          lut[12492] <= 16'd10889;
          lut[12493] <= 16'd10993;
          lut[12494] <= 16'd11096;
          lut[12495] <= 16'd11198;
          lut[12496] <= 16'd11299;
          lut[12497] <= 16'd11399;
          lut[12498] <= 16'd11498;
          lut[12499] <= 16'd11596;
          lut[12500] <= 16'd11693;
          lut[12501] <= 16'd11789;
          lut[12502] <= 16'd11884;
          lut[12503] <= 16'd11978;
          lut[12504] <= 16'd12072;
          lut[12505] <= 16'd12164;
          lut[12506] <= 16'd12255;
          lut[12507] <= 16'd12345;
          lut[12508] <= 16'd12435;
          lut[12509] <= 16'd12523;
          lut[12510] <= 16'd12611;
          lut[12511] <= 16'd12697;
          lut[12512] <= 16'd12783;
          lut[12513] <= 16'd12868;
          lut[12514] <= 16'd12952;
          lut[12515] <= 16'd13035;
          lut[12516] <= 16'd13117;
          lut[12517] <= 16'd13199;
          lut[12518] <= 16'd13280;
          lut[12519] <= 16'd13359;
          lut[12520] <= 16'd13438;
          lut[12521] <= 16'd13516;
          lut[12522] <= 16'd13594;
          lut[12523] <= 16'd13670;
          lut[12524] <= 16'd13746;
          lut[12525] <= 16'd13821;
          lut[12526] <= 16'd13896;
          lut[12527] <= 16'd13969;
          lut[12528] <= 16'd14042;
          lut[12529] <= 16'd14114;
          lut[12530] <= 16'd14185;
          lut[12531] <= 16'd14256;
          lut[12532] <= 16'd14326;
          lut[12533] <= 16'd14395;
          lut[12534] <= 16'd14463;
          lut[12535] <= 16'd14531;
          lut[12536] <= 16'd14598;
          lut[12537] <= 16'd14664;
          lut[12538] <= 16'd14730;
          lut[12539] <= 16'd14795;
          lut[12540] <= 16'd14860;
          lut[12541] <= 16'd14924;
          lut[12542] <= 16'd14987;
          lut[12543] <= 16'd15049;
          lut[12544] <= 0;
          lut[12545] <= 16'd167;
          lut[12546] <= 16'd334;
          lut[12547] <= 16'd501;
          lut[12548] <= 16'd668;
          lut[12549] <= 16'd835;
          lut[12550] <= 16'd1002;
          lut[12551] <= 16'd1168;
          lut[12552] <= 16'd1335;
          lut[12553] <= 16'd1500;
          lut[12554] <= 16'd1666;
          lut[12555] <= 16'd1831;
          lut[12556] <= 16'd1996;
          lut[12557] <= 16'd2161;
          lut[12558] <= 16'd2325;
          lut[12559] <= 16'd2488;
          lut[12560] <= 16'd2652;
          lut[12561] <= 16'd2814;
          lut[12562] <= 16'd2976;
          lut[12563] <= 16'd3138;
          lut[12564] <= 16'd3298;
          lut[12565] <= 16'd3459;
          lut[12566] <= 16'd3618;
          lut[12567] <= 16'd3777;
          lut[12568] <= 16'd3935;
          lut[12569] <= 16'd4092;
          lut[12570] <= 16'd4249;
          lut[12571] <= 16'd4405;
          lut[12572] <= 16'd4560;
          lut[12573] <= 16'd4714;
          lut[12574] <= 16'd4867;
          lut[12575] <= 16'd5020;
          lut[12576] <= 16'd5171;
          lut[12577] <= 16'd5322;
          lut[12578] <= 16'd5471;
          lut[12579] <= 16'd5620;
          lut[12580] <= 16'd5768;
          lut[12581] <= 16'd5915;
          lut[12582] <= 16'd6061;
          lut[12583] <= 16'd6205;
          lut[12584] <= 16'd6349;
          lut[12585] <= 16'd6492;
          lut[12586] <= 16'd6634;
          lut[12587] <= 16'd6774;
          lut[12588] <= 16'd6914;
          lut[12589] <= 16'd7053;
          lut[12590] <= 16'd7190;
          lut[12591] <= 16'd7327;
          lut[12592] <= 16'd7462;
          lut[12593] <= 16'd7596;
          lut[12594] <= 16'd7730;
          lut[12595] <= 16'd7862;
          lut[12596] <= 16'd7993;
          lut[12597] <= 16'd8123;
          lut[12598] <= 16'd8251;
          lut[12599] <= 16'd8379;
          lut[12600] <= 16'd8506;
          lut[12601] <= 16'd8631;
          lut[12602] <= 16'd8756;
          lut[12603] <= 16'd8879;
          lut[12604] <= 16'd9001;
          lut[12605] <= 16'd9122;
          lut[12606] <= 16'd9242;
          lut[12607] <= 16'd9361;
          lut[12608] <= 16'd9479;
          lut[12609] <= 16'd9595;
          lut[12610] <= 16'd9711;
          lut[12611] <= 16'd9825;
          lut[12612] <= 16'd9939;
          lut[12613] <= 16'd10051;
          lut[12614] <= 16'd10162;
          lut[12615] <= 16'd10272;
          lut[12616] <= 16'd10381;
          lut[12617] <= 16'd10489;
          lut[12618] <= 16'd10596;
          lut[12619] <= 16'd10702;
          lut[12620] <= 16'd10807;
          lut[12621] <= 16'd10911;
          lut[12622] <= 16'd11014;
          lut[12623] <= 16'd11116;
          lut[12624] <= 16'd11217;
          lut[12625] <= 16'd11317;
          lut[12626] <= 16'd11415;
          lut[12627] <= 16'd11513;
          lut[12628] <= 16'd11610;
          lut[12629] <= 16'd11706;
          lut[12630] <= 16'd11801;
          lut[12631] <= 16'd11895;
          lut[12632] <= 16'd11988;
          lut[12633] <= 16'd12080;
          lut[12634] <= 16'd12171;
          lut[12635] <= 16'd12261;
          lut[12636] <= 16'd12351;
          lut[12637] <= 16'd12439;
          lut[12638] <= 16'd12527;
          lut[12639] <= 16'd12613;
          lut[12640] <= 16'd12699;
          lut[12641] <= 16'd12784;
          lut[12642] <= 16'd12868;
          lut[12643] <= 16'd12951;
          lut[12644] <= 16'd13033;
          lut[12645] <= 16'd13115;
          lut[12646] <= 16'd13196;
          lut[12647] <= 16'd13275;
          lut[12648] <= 16'd13354;
          lut[12649] <= 16'd13433;
          lut[12650] <= 16'd13510;
          lut[12651] <= 16'd13587;
          lut[12652] <= 16'd13663;
          lut[12653] <= 16'd13738;
          lut[12654] <= 16'd13812;
          lut[12655] <= 16'd13886;
          lut[12656] <= 16'd13959;
          lut[12657] <= 16'd14031;
          lut[12658] <= 16'd14102;
          lut[12659] <= 16'd14173;
          lut[12660] <= 16'd14243;
          lut[12661] <= 16'd14312;
          lut[12662] <= 16'd14381;
          lut[12663] <= 16'd14449;
          lut[12664] <= 16'd14516;
          lut[12665] <= 16'd14582;
          lut[12666] <= 16'd14648;
          lut[12667] <= 16'd14714;
          lut[12668] <= 16'd14778;
          lut[12669] <= 16'd14842;
          lut[12670] <= 16'd14905;
          lut[12671] <= 16'd14968;
          lut[12672] <= 0;
          lut[12673] <= 16'd165;
          lut[12674] <= 16'd331;
          lut[12675] <= 16'd496;
          lut[12676] <= 16'd662;
          lut[12677] <= 16'd827;
          lut[12678] <= 16'd992;
          lut[12679] <= 16'd1157;
          lut[12680] <= 16'd1321;
          lut[12681] <= 16'd1485;
          lut[12682] <= 16'd1649;
          lut[12683] <= 16'd1813;
          lut[12684] <= 16'd1976;
          lut[12685] <= 16'd2139;
          lut[12686] <= 16'd2302;
          lut[12687] <= 16'd2464;
          lut[12688] <= 16'd2625;
          lut[12689] <= 16'd2786;
          lut[12690] <= 16'd2947;
          lut[12691] <= 16'd3107;
          lut[12692] <= 16'd3266;
          lut[12693] <= 16'd3425;
          lut[12694] <= 16'd3583;
          lut[12695] <= 16'd3740;
          lut[12696] <= 16'd3897;
          lut[12697] <= 16'd4053;
          lut[12698] <= 16'd4208;
          lut[12699] <= 16'd4362;
          lut[12700] <= 16'd4516;
          lut[12701] <= 16'd4669;
          lut[12702] <= 16'd4821;
          lut[12703] <= 16'd4972;
          lut[12704] <= 16'd5122;
          lut[12705] <= 16'd5272;
          lut[12706] <= 16'd5420;
          lut[12707] <= 16'd5568;
          lut[12708] <= 16'd5714;
          lut[12709] <= 16'd5860;
          lut[12710] <= 16'd6005;
          lut[12711] <= 16'd6148;
          lut[12712] <= 16'd6291;
          lut[12713] <= 16'd6433;
          lut[12714] <= 16'd6574;
          lut[12715] <= 16'd6713;
          lut[12716] <= 16'd6852;
          lut[12717] <= 16'd6990;
          lut[12718] <= 16'd7126;
          lut[12719] <= 16'd7262;
          lut[12720] <= 16'd7397;
          lut[12721] <= 16'd7530;
          lut[12722] <= 16'd7662;
          lut[12723] <= 16'd7794;
          lut[12724] <= 16'd7924;
          lut[12725] <= 16'd8053;
          lut[12726] <= 16'd8181;
          lut[12727] <= 16'd8308;
          lut[12728] <= 16'd8434;
          lut[12729] <= 16'd8559;
          lut[12730] <= 16'd8683;
          lut[12731] <= 16'd8805;
          lut[12732] <= 16'd8927;
          lut[12733] <= 16'd9048;
          lut[12734] <= 16'd9167;
          lut[12735] <= 16'd9285;
          lut[12736] <= 16'd9403;
          lut[12737] <= 16'd9519;
          lut[12738] <= 16'd9634;
          lut[12739] <= 16'd9748;
          lut[12740] <= 16'd9861;
          lut[12741] <= 16'd9973;
          lut[12742] <= 16'd10084;
          lut[12743] <= 16'd10193;
          lut[12744] <= 16'd10302;
          lut[12745] <= 16'd10410;
          lut[12746] <= 16'd10517;
          lut[12747] <= 16'd10622;
          lut[12748] <= 16'd10727;
          lut[12749] <= 16'd10831;
          lut[12750] <= 16'd10933;
          lut[12751] <= 16'd11035;
          lut[12752] <= 16'd11135;
          lut[12753] <= 16'd11235;
          lut[12754] <= 16'd11334;
          lut[12755] <= 16'd11431;
          lut[12756] <= 16'd11528;
          lut[12757] <= 16'd11624;
          lut[12758] <= 16'd11719;
          lut[12759] <= 16'd11812;
          lut[12760] <= 16'd11905;
          lut[12761] <= 16'd11997;
          lut[12762] <= 16'd12088;
          lut[12763] <= 16'd12179;
          lut[12764] <= 16'd12268;
          lut[12765] <= 16'd12356;
          lut[12766] <= 16'd12444;
          lut[12767] <= 16'd12530;
          lut[12768] <= 16'd12616;
          lut[12769] <= 16'd12701;
          lut[12770] <= 16'd12785;
          lut[12771] <= 16'd12868;
          lut[12772] <= 16'd12950;
          lut[12773] <= 16'd13032;
          lut[12774] <= 16'd13112;
          lut[12775] <= 16'd13192;
          lut[12776] <= 16'd13271;
          lut[12777] <= 16'd13350;
          lut[12778] <= 16'd13427;
          lut[12779] <= 16'd13504;
          lut[12780] <= 16'd13580;
          lut[12781] <= 16'd13655;
          lut[12782] <= 16'd13729;
          lut[12783] <= 16'd13803;
          lut[12784] <= 16'd13876;
          lut[12785] <= 16'd13948;
          lut[12786] <= 16'd14020;
          lut[12787] <= 16'd14091;
          lut[12788] <= 16'd14161;
          lut[12789] <= 16'd14230;
          lut[12790] <= 16'd14299;
          lut[12791] <= 16'd14367;
          lut[12792] <= 16'd14434;
          lut[12793] <= 16'd14501;
          lut[12794] <= 16'd14567;
          lut[12795] <= 16'd14632;
          lut[12796] <= 16'd14697;
          lut[12797] <= 16'd14761;
          lut[12798] <= 16'd14825;
          lut[12799] <= 16'd14888;
          lut[12800] <= 0;
          lut[12801] <= 16'd164;
          lut[12802] <= 16'd328;
          lut[12803] <= 16'd491;
          lut[12804] <= 16'd655;
          lut[12805] <= 16'd819;
          lut[12806] <= 16'd982;
          lut[12807] <= 16'd1145;
          lut[12808] <= 16'd1308;
          lut[12809] <= 16'd1471;
          lut[12810] <= 16'd1633;
          lut[12811] <= 16'd1795;
          lut[12812] <= 16'd1957;
          lut[12813] <= 16'd2118;
          lut[12814] <= 16'd2279;
          lut[12815] <= 16'd2439;
          lut[12816] <= 16'd2599;
          lut[12817] <= 16'd2759;
          lut[12818] <= 16'd2918;
          lut[12819] <= 16'd3076;
          lut[12820] <= 16'd3234;
          lut[12821] <= 16'd3391;
          lut[12822] <= 16'd3548;
          lut[12823] <= 16'd3704;
          lut[12824] <= 16'd3859;
          lut[12825] <= 16'd4014;
          lut[12826] <= 16'd4168;
          lut[12827] <= 16'd4321;
          lut[12828] <= 16'd4473;
          lut[12829] <= 16'd4625;
          lut[12830] <= 16'd4775;
          lut[12831] <= 16'd4925;
          lut[12832] <= 16'd5074;
          lut[12833] <= 16'd5222;
          lut[12834] <= 16'd5370;
          lut[12835] <= 16'd5516;
          lut[12836] <= 16'd5662;
          lut[12837] <= 16'd5806;
          lut[12838] <= 16'd5950;
          lut[12839] <= 16'd6092;
          lut[12840] <= 16'd6234;
          lut[12841] <= 16'd6375;
          lut[12842] <= 16'd6515;
          lut[12843] <= 16'd6654;
          lut[12844] <= 16'd6791;
          lut[12845] <= 16'd6928;
          lut[12846] <= 16'd7064;
          lut[12847] <= 16'd7198;
          lut[12848] <= 16'd7332;
          lut[12849] <= 16'd7465;
          lut[12850] <= 16'd7596;
          lut[12851] <= 16'd7727;
          lut[12852] <= 16'd7856;
          lut[12853] <= 16'd7985;
          lut[12854] <= 16'd8112;
          lut[12855] <= 16'd8239;
          lut[12856] <= 16'd8364;
          lut[12857] <= 16'd8488;
          lut[12858] <= 16'd8611;
          lut[12859] <= 16'd8733;
          lut[12860] <= 16'd8854;
          lut[12861] <= 16'd8974;
          lut[12862] <= 16'd9093;
          lut[12863] <= 16'd9211;
          lut[12864] <= 16'd9328;
          lut[12865] <= 16'd9443;
          lut[12866] <= 16'd9558;
          lut[12867] <= 16'd9672;
          lut[12868] <= 16'd9784;
          lut[12869] <= 16'd9896;
          lut[12870] <= 16'd10006;
          lut[12871] <= 16'd10116;
          lut[12872] <= 16'd10224;
          lut[12873] <= 16'd10331;
          lut[12874] <= 16'd10438;
          lut[12875] <= 16'd10543;
          lut[12876] <= 16'd10647;
          lut[12877] <= 16'd10751;
          lut[12878] <= 16'd10853;
          lut[12879] <= 16'd10955;
          lut[12880] <= 16'd11055;
          lut[12881] <= 16'd11154;
          lut[12882] <= 16'd11253;
          lut[12883] <= 16'd11350;
          lut[12884] <= 16'd11447;
          lut[12885] <= 16'd11542;
          lut[12886] <= 16'd11637;
          lut[12887] <= 16'd11731;
          lut[12888] <= 16'd11824;
          lut[12889] <= 16'd11915;
          lut[12890] <= 16'd12006;
          lut[12891] <= 16'd12097;
          lut[12892] <= 16'd12186;
          lut[12893] <= 16'd12274;
          lut[12894] <= 16'd12361;
          lut[12895] <= 16'd12448;
          lut[12896] <= 16'd12534;
          lut[12897] <= 16'd12618;
          lut[12898] <= 16'd12702;
          lut[12899] <= 16'd12786;
          lut[12900] <= 16'd12868;
          lut[12901] <= 16'd12949;
          lut[12902] <= 16'd13030;
          lut[12903] <= 16'd13110;
          lut[12904] <= 16'd13189;
          lut[12905] <= 16'd13267;
          lut[12906] <= 16'd13345;
          lut[12907] <= 16'd13422;
          lut[12908] <= 16'd13498;
          lut[12909] <= 16'd13573;
          lut[12910] <= 16'd13648;
          lut[12911] <= 16'd13721;
          lut[12912] <= 16'd13794;
          lut[12913] <= 16'd13867;
          lut[12914] <= 16'd13938;
          lut[12915] <= 16'd14009;
          lut[12916] <= 16'd14079;
          lut[12917] <= 16'd14149;
          lut[12918] <= 16'd14218;
          lut[12919] <= 16'd14286;
          lut[12920] <= 16'd14353;
          lut[12921] <= 16'd14420;
          lut[12922] <= 16'd14486;
          lut[12923] <= 16'd14552;
          lut[12924] <= 16'd14617;
          lut[12925] <= 16'd14681;
          lut[12926] <= 16'd14745;
          lut[12927] <= 16'd14808;
          lut[12928] <= 0;
          lut[12929] <= 16'd162;
          lut[12930] <= 16'd324;
          lut[12931] <= 16'd487;
          lut[12932] <= 16'd649;
          lut[12933] <= 16'd810;
          lut[12934] <= 16'd972;
          lut[12935] <= 16'd1134;
          lut[12936] <= 16'd1295;
          lut[12937] <= 16'd1456;
          lut[12938] <= 16'd1617;
          lut[12939] <= 16'd1777;
          lut[12940] <= 16'd1938;
          lut[12941] <= 16'd2097;
          lut[12942] <= 16'd2257;
          lut[12943] <= 16'd2416;
          lut[12944] <= 16'd2574;
          lut[12945] <= 16'd2732;
          lut[12946] <= 16'd2890;
          lut[12947] <= 16'd3047;
          lut[12948] <= 16'd3203;
          lut[12949] <= 16'd3359;
          lut[12950] <= 16'd3514;
          lut[12951] <= 16'd3668;
          lut[12952] <= 16'd3822;
          lut[12953] <= 16'd3976;
          lut[12954] <= 16'd4128;
          lut[12955] <= 16'd4280;
          lut[12956] <= 16'd4431;
          lut[12957] <= 16'd4581;
          lut[12958] <= 16'd4731;
          lut[12959] <= 16'd4879;
          lut[12960] <= 16'd5027;
          lut[12961] <= 16'd5174;
          lut[12962] <= 16'd5320;
          lut[12963] <= 16'd5465;
          lut[12964] <= 16'd5610;
          lut[12965] <= 16'd5753;
          lut[12966] <= 16'd5896;
          lut[12967] <= 16'd6038;
          lut[12968] <= 16'd6178;
          lut[12969] <= 16'd6318;
          lut[12970] <= 16'd6457;
          lut[12971] <= 16'd6595;
          lut[12972] <= 16'd6731;
          lut[12973] <= 16'd6867;
          lut[12974] <= 16'd7002;
          lut[12975] <= 16'd7136;
          lut[12976] <= 16'd7269;
          lut[12977] <= 16'd7401;
          lut[12978] <= 16'd7531;
          lut[12979] <= 16'd7661;
          lut[12980] <= 16'd7790;
          lut[12981] <= 16'd7918;
          lut[12982] <= 16'd8044;
          lut[12983] <= 16'd8170;
          lut[12984] <= 16'd8295;
          lut[12985] <= 16'd8418;
          lut[12986] <= 16'd8541;
          lut[12987] <= 16'd8662;
          lut[12988] <= 16'd8782;
          lut[12989] <= 16'd8902;
          lut[12990] <= 16'd9020;
          lut[12991] <= 16'd9138;
          lut[12992] <= 16'd9254;
          lut[12993] <= 16'd9369;
          lut[12994] <= 16'd9483;
          lut[12995] <= 16'd9596;
          lut[12996] <= 16'd9708;
          lut[12997] <= 16'd9820;
          lut[12998] <= 16'd9930;
          lut[12999] <= 16'd10039;
          lut[13000] <= 16'd10147;
          lut[13001] <= 16'd10254;
          lut[13002] <= 16'd10360;
          lut[13003] <= 16'd10465;
          lut[13004] <= 16'd10569;
          lut[13005] <= 16'd10672;
          lut[13006] <= 16'd10774;
          lut[13007] <= 16'd10875;
          lut[13008] <= 16'd10976;
          lut[13009] <= 16'd11075;
          lut[13010] <= 16'd11173;
          lut[13011] <= 16'd11270;
          lut[13012] <= 16'd11367;
          lut[13013] <= 16'd11462;
          lut[13014] <= 16'd11557;
          lut[13015] <= 16'd11650;
          lut[13016] <= 16'd11743;
          lut[13017] <= 16'd11835;
          lut[13018] <= 16'd11925;
          lut[13019] <= 16'd12015;
          lut[13020] <= 16'd12104;
          lut[13021] <= 16'd12193;
          lut[13022] <= 16'd12280;
          lut[13023] <= 16'd12367;
          lut[13024] <= 16'd12452;
          lut[13025] <= 16'd12537;
          lut[13026] <= 16'd12621;
          lut[13027] <= 16'd12704;
          lut[13028] <= 16'd12786;
          lut[13029] <= 16'd12868;
          lut[13030] <= 16'd12949;
          lut[13031] <= 16'd13029;
          lut[13032] <= 16'd13108;
          lut[13033] <= 16'd13186;
          lut[13034] <= 16'd13264;
          lut[13035] <= 16'd13340;
          lut[13036] <= 16'd13417;
          lut[13037] <= 16'd13492;
          lut[13038] <= 16'd13566;
          lut[13039] <= 16'd13640;
          lut[13040] <= 16'd13713;
          lut[13041] <= 16'd13786;
          lut[13042] <= 16'd13857;
          lut[13043] <= 16'd13928;
          lut[13044] <= 16'd13999;
          lut[13045] <= 16'd14068;
          lut[13046] <= 16'd14137;
          lut[13047] <= 16'd14205;
          lut[13048] <= 16'd14273;
          lut[13049] <= 16'd14340;
          lut[13050] <= 16'd14406;
          lut[13051] <= 16'd14472;
          lut[13052] <= 16'd14537;
          lut[13053] <= 16'd14601;
          lut[13054] <= 16'd14665;
          lut[13055] <= 16'd14728;
          lut[13056] <= 0;
          lut[13057] <= 16'd161;
          lut[13058] <= 16'd321;
          lut[13059] <= 16'd482;
          lut[13060] <= 16'd642;
          lut[13061] <= 16'd802;
          lut[13062] <= 16'd963;
          lut[13063] <= 16'd1123;
          lut[13064] <= 16'd1282;
          lut[13065] <= 16'd1442;
          lut[13066] <= 16'd1601;
          lut[13067] <= 16'd1760;
          lut[13068] <= 16'd1919;
          lut[13069] <= 16'd2077;
          lut[13070] <= 16'd2235;
          lut[13071] <= 16'd2392;
          lut[13072] <= 16'd2549;
          lut[13073] <= 16'd2706;
          lut[13074] <= 16'd2862;
          lut[13075] <= 16'd3017;
          lut[13076] <= 16'd3172;
          lut[13077] <= 16'd3327;
          lut[13078] <= 16'd3480;
          lut[13079] <= 16'd3634;
          lut[13080] <= 16'd3786;
          lut[13081] <= 16'd3938;
          lut[13082] <= 16'd4089;
          lut[13083] <= 16'd4240;
          lut[13084] <= 16'd4389;
          lut[13085] <= 16'd4538;
          lut[13086] <= 16'd4687;
          lut[13087] <= 16'd4834;
          lut[13088] <= 16'd4981;
          lut[13089] <= 16'd5127;
          lut[13090] <= 16'd5272;
          lut[13091] <= 16'd5416;
          lut[13092] <= 16'd5559;
          lut[13093] <= 16'd5701;
          lut[13094] <= 16'd5843;
          lut[13095] <= 16'd5983;
          lut[13096] <= 16'd6123;
          lut[13097] <= 16'd6262;
          lut[13098] <= 16'd6400;
          lut[13099] <= 16'd6537;
          lut[13100] <= 16'd6672;
          lut[13101] <= 16'd6807;
          lut[13102] <= 16'd6941;
          lut[13103] <= 16'd7074;
          lut[13104] <= 16'd7206;
          lut[13105] <= 16'd7337;
          lut[13106] <= 16'd7467;
          lut[13107] <= 16'd7596;
          lut[13108] <= 16'd7724;
          lut[13109] <= 16'd7851;
          lut[13110] <= 16'd7977;
          lut[13111] <= 16'd8102;
          lut[13112] <= 16'd8226;
          lut[13113] <= 16'd8349;
          lut[13114] <= 16'd8471;
          lut[13115] <= 16'd8592;
          lut[13116] <= 16'd8712;
          lut[13117] <= 16'd8831;
          lut[13118] <= 16'd8948;
          lut[13119] <= 16'd9065;
          lut[13120] <= 16'd9181;
          lut[13121] <= 16'd9296;
          lut[13122] <= 16'd9409;
          lut[13123] <= 16'd9522;
          lut[13124] <= 16'd9634;
          lut[13125] <= 16'd9745;
          lut[13126] <= 16'd9854;
          lut[13127] <= 16'd9963;
          lut[13128] <= 16'd10071;
          lut[13129] <= 16'd10177;
          lut[13130] <= 16'd10283;
          lut[13131] <= 16'd10388;
          lut[13132] <= 16'd10492;
          lut[13133] <= 16'd10594;
          lut[13134] <= 16'd10696;
          lut[13135] <= 16'd10797;
          lut[13136] <= 16'd10897;
          lut[13137] <= 16'd10996;
          lut[13138] <= 16'd11094;
          lut[13139] <= 16'd11191;
          lut[13140] <= 16'd11287;
          lut[13141] <= 16'd11383;
          lut[13142] <= 16'd11477;
          lut[13143] <= 16'd11570;
          lut[13144] <= 16'd11663;
          lut[13145] <= 16'd11755;
          lut[13146] <= 16'd11845;
          lut[13147] <= 16'd11935;
          lut[13148] <= 16'd12024;
          lut[13149] <= 16'd12112;
          lut[13150] <= 16'd12200;
          lut[13151] <= 16'd12286;
          lut[13152] <= 16'd12372;
          lut[13153] <= 16'd12456;
          lut[13154] <= 16'd12540;
          lut[13155] <= 16'd12623;
          lut[13156] <= 16'd12706;
          lut[13157] <= 16'd12787;
          lut[13158] <= 16'd12868;
          lut[13159] <= 16'd12948;
          lut[13160] <= 16'd13027;
          lut[13161] <= 16'd13105;
          lut[13162] <= 16'd13183;
          lut[13163] <= 16'd13260;
          lut[13164] <= 16'd13336;
          lut[13165] <= 16'd13411;
          lut[13166] <= 16'd13486;
          lut[13167] <= 16'd13560;
          lut[13168] <= 16'd13633;
          lut[13169] <= 16'd13705;
          lut[13170] <= 16'd13777;
          lut[13171] <= 16'd13848;
          lut[13172] <= 16'd13919;
          lut[13173] <= 16'd13988;
          lut[13174] <= 16'd14057;
          lut[13175] <= 16'd14126;
          lut[13176] <= 16'd14193;
          lut[13177] <= 16'd14261;
          lut[13178] <= 16'd14327;
          lut[13179] <= 16'd14393;
          lut[13180] <= 16'd14458;
          lut[13181] <= 16'd14522;
          lut[13182] <= 16'd14586;
          lut[13183] <= 16'd14650;
          lut[13184] <= 0;
          lut[13185] <= 16'd159;
          lut[13186] <= 16'd318;
          lut[13187] <= 16'd477;
          lut[13188] <= 16'd636;
          lut[13189] <= 16'd795;
          lut[13190] <= 16'd953;
          lut[13191] <= 16'd1112;
          lut[13192] <= 16'd1270;
          lut[13193] <= 16'd1428;
          lut[13194] <= 16'd1586;
          lut[13195] <= 16'd1743;
          lut[13196] <= 16'd1900;
          lut[13197] <= 16'd2057;
          lut[13198] <= 16'd2213;
          lut[13199] <= 16'd2369;
          lut[13200] <= 16'd2525;
          lut[13201] <= 16'd2680;
          lut[13202] <= 16'd2835;
          lut[13203] <= 16'd2989;
          lut[13204] <= 16'd3142;
          lut[13205] <= 16'd3295;
          lut[13206] <= 16'd3448;
          lut[13207] <= 16'd3600;
          lut[13208] <= 16'd3751;
          lut[13209] <= 16'd3901;
          lut[13210] <= 16'd4051;
          lut[13211] <= 16'd4200;
          lut[13212] <= 16'd4349;
          lut[13213] <= 16'd4497;
          lut[13214] <= 16'd4644;
          lut[13215] <= 16'd4790;
          lut[13216] <= 16'd4935;
          lut[13217] <= 16'd5080;
          lut[13218] <= 16'd5224;
          lut[13219] <= 16'd5367;
          lut[13220] <= 16'd5509;
          lut[13221] <= 16'd5650;
          lut[13222] <= 16'd5791;
          lut[13223] <= 16'd5930;
          lut[13224] <= 16'd6069;
          lut[13225] <= 16'd6207;
          lut[13226] <= 16'd6344;
          lut[13227] <= 16'd6480;
          lut[13228] <= 16'd6615;
          lut[13229] <= 16'd6749;
          lut[13230] <= 16'd6882;
          lut[13231] <= 16'd7014;
          lut[13232] <= 16'd7145;
          lut[13233] <= 16'd7275;
          lut[13234] <= 16'd7404;
          lut[13235] <= 16'd7533;
          lut[13236] <= 16'd7660;
          lut[13237] <= 16'd7786;
          lut[13238] <= 16'd7911;
          lut[13239] <= 16'd8036;
          lut[13240] <= 16'd8159;
          lut[13241] <= 16'd8281;
          lut[13242] <= 16'd8403;
          lut[13243] <= 16'd8523;
          lut[13244] <= 16'd8642;
          lut[13245] <= 16'd8760;
          lut[13246] <= 16'd8878;
          lut[13247] <= 16'd8994;
          lut[13248] <= 16'd9109;
          lut[13249] <= 16'd9223;
          lut[13250] <= 16'd9337;
          lut[13251] <= 16'd9449;
          lut[13252] <= 16'd9560;
          lut[13253] <= 16'd9670;
          lut[13254] <= 16'd9780;
          lut[13255] <= 16'd9888;
          lut[13256] <= 16'd9995;
          lut[13257] <= 16'd10102;
          lut[13258] <= 16'd10207;
          lut[13259] <= 16'd10312;
          lut[13260] <= 16'd10415;
          lut[13261] <= 16'd10518;
          lut[13262] <= 16'd10619;
          lut[13263] <= 16'd10720;
          lut[13264] <= 16'd10820;
          lut[13265] <= 16'd10918;
          lut[13266] <= 16'd11016;
          lut[13267] <= 16'd11113;
          lut[13268] <= 16'd11209;
          lut[13269] <= 16'd11304;
          lut[13270] <= 16'd11398;
          lut[13271] <= 16'd11492;
          lut[13272] <= 16'd11584;
          lut[13273] <= 16'd11675;
          lut[13274] <= 16'd11766;
          lut[13275] <= 16'd11856;
          lut[13276] <= 16'd11945;
          lut[13277] <= 16'd12033;
          lut[13278] <= 16'd12120;
          lut[13279] <= 16'd12206;
          lut[13280] <= 16'd12292;
          lut[13281] <= 16'd12377;
          lut[13282] <= 16'd12460;
          lut[13283] <= 16'd12544;
          lut[13284] <= 16'd12626;
          lut[13285] <= 16'd12707;
          lut[13286] <= 16'd12788;
          lut[13287] <= 16'd12868;
          lut[13288] <= 16'd12947;
          lut[13289] <= 16'd13025;
          lut[13290] <= 16'd13103;
          lut[13291] <= 16'd13180;
          lut[13292] <= 16'd13256;
          lut[13293] <= 16'd13332;
          lut[13294] <= 16'd13406;
          lut[13295] <= 16'd13480;
          lut[13296] <= 16'd13553;
          lut[13297] <= 16'd13626;
          lut[13298] <= 16'd13698;
          lut[13299] <= 16'd13769;
          lut[13300] <= 16'd13839;
          lut[13301] <= 16'd13909;
          lut[13302] <= 16'd13978;
          lut[13303] <= 16'd14047;
          lut[13304] <= 16'd14115;
          lut[13305] <= 16'd14182;
          lut[13306] <= 16'd14248;
          lut[13307] <= 16'd14314;
          lut[13308] <= 16'd14379;
          lut[13309] <= 16'd14444;
          lut[13310] <= 16'd14508;
          lut[13311] <= 16'd14571;
          lut[13312] <= 0;
          lut[13313] <= 16'd158;
          lut[13314] <= 16'd315;
          lut[13315] <= 16'd472;
          lut[13316] <= 16'd630;
          lut[13317] <= 16'd787;
          lut[13318] <= 16'd944;
          lut[13319] <= 16'd1101;
          lut[13320] <= 16'd1258;
          lut[13321] <= 16'd1414;
          lut[13322] <= 16'd1571;
          lut[13323] <= 16'd1727;
          lut[13324] <= 16'd1882;
          lut[13325] <= 16'd2037;
          lut[13326] <= 16'd2192;
          lut[13327] <= 16'd2347;
          lut[13328] <= 16'd2501;
          lut[13329] <= 16'd2655;
          lut[13330] <= 16'd2808;
          lut[13331] <= 16'd2961;
          lut[13332] <= 16'd3113;
          lut[13333] <= 16'd3264;
          lut[13334] <= 16'd3415;
          lut[13335] <= 16'd3566;
          lut[13336] <= 16'd3716;
          lut[13337] <= 16'd3865;
          lut[13338] <= 16'd4014;
          lut[13339] <= 16'd4162;
          lut[13340] <= 16'd4309;
          lut[13341] <= 16'd4455;
          lut[13342] <= 16'd4601;
          lut[13343] <= 16'd4746;
          lut[13344] <= 16'd4891;
          lut[13345] <= 16'd5034;
          lut[13346] <= 16'd5177;
          lut[13347] <= 16'd5319;
          lut[13348] <= 16'd5460;
          lut[13349] <= 16'd5600;
          lut[13350] <= 16'd5740;
          lut[13351] <= 16'd5878;
          lut[13352] <= 16'd6016;
          lut[13353] <= 16'd6153;
          lut[13354] <= 16'd6288;
          lut[13355] <= 16'd6423;
          lut[13356] <= 16'd6558;
          lut[13357] <= 16'd6691;
          lut[13358] <= 16'd6823;
          lut[13359] <= 16'd6954;
          lut[13360] <= 16'd7085;
          lut[13361] <= 16'd7214;
          lut[13362] <= 16'd7342;
          lut[13363] <= 16'd7470;
          lut[13364] <= 16'd7596;
          lut[13365] <= 16'd7722;
          lut[13366] <= 16'd7847;
          lut[13367] <= 16'd7970;
          lut[13368] <= 16'd8093;
          lut[13369] <= 16'd8214;
          lut[13370] <= 16'd8335;
          lut[13371] <= 16'd8455;
          lut[13372] <= 16'd8573;
          lut[13373] <= 16'd8691;
          lut[13374] <= 16'd8808;
          lut[13375] <= 16'd8924;
          lut[13376] <= 16'd9038;
          lut[13377] <= 16'd9152;
          lut[13378] <= 16'd9265;
          lut[13379] <= 16'd9377;
          lut[13380] <= 16'd9488;
          lut[13381] <= 16'd9597;
          lut[13382] <= 16'd9706;
          lut[13383] <= 16'd9814;
          lut[13384] <= 16'd9921;
          lut[13385] <= 16'd10027;
          lut[13386] <= 16'd10132;
          lut[13387] <= 16'd10236;
          lut[13388] <= 16'd10340;
          lut[13389] <= 16'd10442;
          lut[13390] <= 16'd10543;
          lut[13391] <= 16'd10643;
          lut[13392] <= 16'd10743;
          lut[13393] <= 16'd10841;
          lut[13394] <= 16'd10939;
          lut[13395] <= 16'd11036;
          lut[13396] <= 16'd11132;
          lut[13397] <= 16'd11226;
          lut[13398] <= 16'd11320;
          lut[13399] <= 16'd11414;
          lut[13400] <= 16'd11506;
          lut[13401] <= 16'd11597;
          lut[13402] <= 16'd11688;
          lut[13403] <= 16'd11777;
          lut[13404] <= 16'd11866;
          lut[13405] <= 16'd11954;
          lut[13406] <= 16'd12041;
          lut[13407] <= 16'd12127;
          lut[13408] <= 16'd12213;
          lut[13409] <= 16'd12298;
          lut[13410] <= 16'd12381;
          lut[13411] <= 16'd12464;
          lut[13412] <= 16'd12547;
          lut[13413] <= 16'd12628;
          lut[13414] <= 16'd12709;
          lut[13415] <= 16'd12789;
          lut[13416] <= 16'd12868;
          lut[13417] <= 16'd12946;
          lut[13418] <= 16'd13024;
          lut[13419] <= 16'd13101;
          lut[13420] <= 16'd13177;
          lut[13421] <= 16'd13252;
          lut[13422] <= 16'd13327;
          lut[13423] <= 16'd13401;
          lut[13424] <= 16'd13475;
          lut[13425] <= 16'd13547;
          lut[13426] <= 16'd13619;
          lut[13427] <= 16'd13690;
          lut[13428] <= 16'd13761;
          lut[13429] <= 16'd13831;
          lut[13430] <= 16'd13900;
          lut[13431] <= 16'd13968;
          lut[13432] <= 16'd14036;
          lut[13433] <= 16'd14104;
          lut[13434] <= 16'd14170;
          lut[13435] <= 16'd14236;
          lut[13436] <= 16'd14301;
          lut[13437] <= 16'd14366;
          lut[13438] <= 16'd14430;
          lut[13439] <= 16'd14494;
          lut[13440] <= 0;
          lut[13441] <= 16'd156;
          lut[13442] <= 16'd312;
          lut[13443] <= 16'd468;
          lut[13444] <= 16'd624;
          lut[13445] <= 16'd780;
          lut[13446] <= 16'd935;
          lut[13447] <= 16'd1091;
          lut[13448] <= 16'd1246;
          lut[13449] <= 16'd1401;
          lut[13450] <= 16'd1556;
          lut[13451] <= 16'd1710;
          lut[13452] <= 16'd1864;
          lut[13453] <= 16'd2018;
          lut[13454] <= 16'd2172;
          lut[13455] <= 16'd2325;
          lut[13456] <= 16'd2478;
          lut[13457] <= 16'd2630;
          lut[13458] <= 16'd2782;
          lut[13459] <= 16'd2933;
          lut[13460] <= 16'd3084;
          lut[13461] <= 16'd3234;
          lut[13462] <= 16'd3384;
          lut[13463] <= 16'd3533;
          lut[13464] <= 16'd3682;
          lut[13465] <= 16'd3830;
          lut[13466] <= 16'd3977;
          lut[13467] <= 16'd4124;
          lut[13468] <= 16'd4270;
          lut[13469] <= 16'd4415;
          lut[13470] <= 16'd4560;
          lut[13471] <= 16'd4704;
          lut[13472] <= 16'd4847;
          lut[13473] <= 16'd4989;
          lut[13474] <= 16'd5131;
          lut[13475] <= 16'd5272;
          lut[13476] <= 16'd5412;
          lut[13477] <= 16'd5551;
          lut[13478] <= 16'd5689;
          lut[13479] <= 16'd5827;
          lut[13480] <= 16'd5963;
          lut[13481] <= 16'd6099;
          lut[13482] <= 16'd6234;
          lut[13483] <= 16'd6368;
          lut[13484] <= 16'd6501;
          lut[13485] <= 16'd6634;
          lut[13486] <= 16'd6765;
          lut[13487] <= 16'd6896;
          lut[13488] <= 16'd7025;
          lut[13489] <= 16'd7154;
          lut[13490] <= 16'd7281;
          lut[13491] <= 16'd7408;
          lut[13492] <= 16'd7534;
          lut[13493] <= 16'd7659;
          lut[13494] <= 16'd7783;
          lut[13495] <= 16'd7905;
          lut[13496] <= 16'd8027;
          lut[13497] <= 16'd8148;
          lut[13498] <= 16'd8269;
          lut[13499] <= 16'd8388;
          lut[13500] <= 16'd8506;
          lut[13501] <= 16'd8623;
          lut[13502] <= 16'd8739;
          lut[13503] <= 16'd8854;
          lut[13504] <= 16'd8968;
          lut[13505] <= 16'd9082;
          lut[13506] <= 16'd9194;
          lut[13507] <= 16'd9305;
          lut[13508] <= 16'd9416;
          lut[13509] <= 16'd9525;
          lut[13510] <= 16'd9634;
          lut[13511] <= 16'd9741;
          lut[13512] <= 16'd9848;
          lut[13513] <= 16'd9954;
          lut[13514] <= 16'd10058;
          lut[13515] <= 16'd10162;
          lut[13516] <= 16'd10265;
          lut[13517] <= 16'd10367;
          lut[13518] <= 16'd10468;
          lut[13519] <= 16'd10568;
          lut[13520] <= 16'd10667;
          lut[13521] <= 16'd10766;
          lut[13522] <= 16'd10863;
          lut[13523] <= 16'd10959;
          lut[13524] <= 16'd11055;
          lut[13525] <= 16'd11150;
          lut[13526] <= 16'd11243;
          lut[13527] <= 16'd11336;
          lut[13528] <= 16'd11429;
          lut[13529] <= 16'd11520;
          lut[13530] <= 16'd11610;
          lut[13531] <= 16'd11700;
          lut[13532] <= 16'd11788;
          lut[13533] <= 16'd11876;
          lut[13534] <= 16'd11963;
          lut[13535] <= 16'd12049;
          lut[13536] <= 16'd12135;
          lut[13537] <= 16'd12219;
          lut[13538] <= 16'd12303;
          lut[13539] <= 16'd12386;
          lut[13540] <= 16'd12468;
          lut[13541] <= 16'd12550;
          lut[13542] <= 16'd12631;
          lut[13543] <= 16'd12710;
          lut[13544] <= 16'd12790;
          lut[13545] <= 16'd12868;
          lut[13546] <= 16'd12946;
          lut[13547] <= 16'd13023;
          lut[13548] <= 16'd13099;
          lut[13549] <= 16'd13174;
          lut[13550] <= 16'd13249;
          lut[13551] <= 16'd13323;
          lut[13552] <= 16'd13396;
          lut[13553] <= 16'd13469;
          lut[13554] <= 16'd13541;
          lut[13555] <= 16'd13612;
          lut[13556] <= 16'd13683;
          lut[13557] <= 16'd13753;
          lut[13558] <= 16'd13822;
          lut[13559] <= 16'd13891;
          lut[13560] <= 16'd13959;
          lut[13561] <= 16'd14026;
          lut[13562] <= 16'd14093;
          lut[13563] <= 16'd14159;
          lut[13564] <= 16'd14224;
          lut[13565] <= 16'd14289;
          lut[13566] <= 16'd14353;
          lut[13567] <= 16'd14417;
          lut[13568] <= 0;
          lut[13569] <= 16'd155;
          lut[13570] <= 16'd309;
          lut[13571] <= 16'd464;
          lut[13572] <= 16'd618;
          lut[13573] <= 16'd772;
          lut[13574] <= 16'd926;
          lut[13575] <= 16'd1080;
          lut[13576] <= 16'd1234;
          lut[13577] <= 16'd1388;
          lut[13578] <= 16'd1541;
          lut[13579] <= 16'd1694;
          lut[13580] <= 16'd1847;
          lut[13581] <= 16'd1999;
          lut[13582] <= 16'd2151;
          lut[13583] <= 16'd2303;
          lut[13584] <= 16'd2455;
          lut[13585] <= 16'd2605;
          lut[13586] <= 16'd2756;
          lut[13587] <= 16'd2906;
          lut[13588] <= 16'd3055;
          lut[13589] <= 16'd3204;
          lut[13590] <= 16'd3353;
          lut[13591] <= 16'd3501;
          lut[13592] <= 16'd3648;
          lut[13593] <= 16'd3795;
          lut[13594] <= 16'd3941;
          lut[13595] <= 16'd4086;
          lut[13596] <= 16'd4231;
          lut[13597] <= 16'd4375;
          lut[13598] <= 16'd4519;
          lut[13599] <= 16'd4662;
          lut[13600] <= 16'd4804;
          lut[13601] <= 16'd4945;
          lut[13602] <= 16'd5085;
          lut[13603] <= 16'd5225;
          lut[13604] <= 16'd5364;
          lut[13605] <= 16'd5502;
          lut[13606] <= 16'd5640;
          lut[13607] <= 16'd5776;
          lut[13608] <= 16'd5912;
          lut[13609] <= 16'd6047;
          lut[13610] <= 16'd6181;
          lut[13611] <= 16'd6314;
          lut[13612] <= 16'd6446;
          lut[13613] <= 16'd6578;
          lut[13614] <= 16'd6708;
          lut[13615] <= 16'd6838;
          lut[13616] <= 16'd6967;
          lut[13617] <= 16'd7094;
          lut[13618] <= 16'd7221;
          lut[13619] <= 16'd7347;
          lut[13620] <= 16'd7472;
          lut[13621] <= 16'd7596;
          lut[13622] <= 16'd7720;
          lut[13623] <= 16'd7842;
          lut[13624] <= 16'd7963;
          lut[13625] <= 16'd8084;
          lut[13626] <= 16'd8203;
          lut[13627] <= 16'd8321;
          lut[13628] <= 16'd8439;
          lut[13629] <= 16'd8556;
          lut[13630] <= 16'd8671;
          lut[13631] <= 16'd8786;
          lut[13632] <= 16'd8900;
          lut[13633] <= 16'd9012;
          lut[13634] <= 16'd9124;
          lut[13635] <= 16'd9235;
          lut[13636] <= 16'd9345;
          lut[13637] <= 16'd9454;
          lut[13638] <= 16'd9562;
          lut[13639] <= 16'd9669;
          lut[13640] <= 16'd9776;
          lut[13641] <= 16'd9881;
          lut[13642] <= 16'd9985;
          lut[13643] <= 16'd10089;
          lut[13644] <= 16'd10191;
          lut[13645] <= 16'd10293;
          lut[13646] <= 16'd10394;
          lut[13647] <= 16'd10494;
          lut[13648] <= 16'd10592;
          lut[13649] <= 16'd10691;
          lut[13650] <= 16'd10788;
          lut[13651] <= 16'd10884;
          lut[13652] <= 16'd10979;
          lut[13653] <= 16'd11074;
          lut[13654] <= 16'd11167;
          lut[13655] <= 16'd11260;
          lut[13656] <= 16'd11352;
          lut[13657] <= 16'd11443;
          lut[13658] <= 16'd11533;
          lut[13659] <= 16'd11623;
          lut[13660] <= 16'd11711;
          lut[13661] <= 16'd11799;
          lut[13662] <= 16'd11886;
          lut[13663] <= 16'd11972;
          lut[13664] <= 16'd12058;
          lut[13665] <= 16'd12142;
          lut[13666] <= 16'd12226;
          lut[13667] <= 16'd12309;
          lut[13668] <= 16'd12391;
          lut[13669] <= 16'd12472;
          lut[13670] <= 16'd12553;
          lut[13671] <= 16'd12633;
          lut[13672] <= 16'd12712;
          lut[13673] <= 16'd12790;
          lut[13674] <= 16'd12868;
          lut[13675] <= 16'd12945;
          lut[13676] <= 16'd13021;
          lut[13677] <= 16'd13097;
          lut[13678] <= 16'd13171;
          lut[13679] <= 16'd13245;
          lut[13680] <= 16'd13319;
          lut[13681] <= 16'd13391;
          lut[13682] <= 16'd13463;
          lut[13683] <= 16'd13535;
          lut[13684] <= 16'd13605;
          lut[13685] <= 16'd13675;
          lut[13686] <= 16'd13745;
          lut[13687] <= 16'd13814;
          lut[13688] <= 16'd13882;
          lut[13689] <= 16'd13949;
          lut[13690] <= 16'd14016;
          lut[13691] <= 16'd14082;
          lut[13692] <= 16'd14148;
          lut[13693] <= 16'd14213;
          lut[13694] <= 16'd14277;
          lut[13695] <= 16'd14341;
          lut[13696] <= 0;
          lut[13697] <= 16'd153;
          lut[13698] <= 16'd306;
          lut[13699] <= 16'd459;
          lut[13700] <= 16'd612;
          lut[13701] <= 16'd765;
          lut[13702] <= 16'd918;
          lut[13703] <= 16'd1070;
          lut[13704] <= 16'd1223;
          lut[13705] <= 16'd1375;
          lut[13706] <= 16'd1527;
          lut[13707] <= 16'd1678;
          lut[13708] <= 16'd1830;
          lut[13709] <= 16'd1981;
          lut[13710] <= 16'd2132;
          lut[13711] <= 16'd2282;
          lut[13712] <= 16'd2432;
          lut[13713] <= 16'd2581;
          lut[13714] <= 16'd2731;
          lut[13715] <= 16'd2879;
          lut[13716] <= 16'd3027;
          lut[13717] <= 16'd3175;
          lut[13718] <= 16'd3322;
          lut[13719] <= 16'd3469;
          lut[13720] <= 16'd3615;
          lut[13721] <= 16'd3761;
          lut[13722] <= 16'd3905;
          lut[13723] <= 16'd4050;
          lut[13724] <= 16'd4193;
          lut[13725] <= 16'd4336;
          lut[13726] <= 16'd4479;
          lut[13727] <= 16'd4620;
          lut[13728] <= 16'd4761;
          lut[13729] <= 16'd4901;
          lut[13730] <= 16'd5041;
          lut[13731] <= 16'd5180;
          lut[13732] <= 16'd5317;
          lut[13733] <= 16'd5455;
          lut[13734] <= 16'd5591;
          lut[13735] <= 16'd5727;
          lut[13736] <= 16'd5861;
          lut[13737] <= 16'd5995;
          lut[13738] <= 16'd6128;
          lut[13739] <= 16'd6261;
          lut[13740] <= 16'd6392;
          lut[13741] <= 16'd6523;
          lut[13742] <= 16'd6652;
          lut[13743] <= 16'd6781;
          lut[13744] <= 16'd6909;
          lut[13745] <= 16'd7036;
          lut[13746] <= 16'd7162;
          lut[13747] <= 16'd7287;
          lut[13748] <= 16'd7412;
          lut[13749] <= 16'd7535;
          lut[13750] <= 16'd7658;
          lut[13751] <= 16'd7779;
          lut[13752] <= 16'd7900;
          lut[13753] <= 16'd8020;
          lut[13754] <= 16'd8138;
          lut[13755] <= 16'd8256;
          lut[13756] <= 16'd8373;
          lut[13757] <= 16'd8489;
          lut[13758] <= 16'd8604;
          lut[13759] <= 16'd8718;
          lut[13760] <= 16'd8832;
          lut[13761] <= 16'd8944;
          lut[13762] <= 16'd9055;
          lut[13763] <= 16'd9166;
          lut[13764] <= 16'd9275;
          lut[13765] <= 16'd9384;
          lut[13766] <= 16'd9492;
          lut[13767] <= 16'd9598;
          lut[13768] <= 16'd9704;
          lut[13769] <= 16'd9809;
          lut[13770] <= 16'd9913;
          lut[13771] <= 16'd10016;
          lut[13772] <= 16'd10119;
          lut[13773] <= 16'd10220;
          lut[13774] <= 16'd10320;
          lut[13775] <= 16'd10420;
          lut[13776] <= 16'd10519;
          lut[13777] <= 16'd10616;
          lut[13778] <= 16'd10713;
          lut[13779] <= 16'd10809;
          lut[13780] <= 16'd10904;
          lut[13781] <= 16'd10999;
          lut[13782] <= 16'd11092;
          lut[13783] <= 16'd11185;
          lut[13784] <= 16'd11277;
          lut[13785] <= 16'd11368;
          lut[13786] <= 16'd11458;
          lut[13787] <= 16'd11547;
          lut[13788] <= 16'd11635;
          lut[13789] <= 16'd11723;
          lut[13790] <= 16'd11810;
          lut[13791] <= 16'd11896;
          lut[13792] <= 16'd11981;
          lut[13793] <= 16'd12065;
          lut[13794] <= 16'd12149;
          lut[13795] <= 16'd12232;
          lut[13796] <= 16'd12314;
          lut[13797] <= 16'd12395;
          lut[13798] <= 16'd12476;
          lut[13799] <= 16'd12556;
          lut[13800] <= 16'd12635;
          lut[13801] <= 16'd12713;
          lut[13802] <= 16'd12791;
          lut[13803] <= 16'd12868;
          lut[13804] <= 16'd12944;
          lut[13805] <= 16'd13020;
          lut[13806] <= 16'd13094;
          lut[13807] <= 16'd13169;
          lut[13808] <= 16'd13242;
          lut[13809] <= 16'd13315;
          lut[13810] <= 16'd13387;
          lut[13811] <= 16'd13458;
          lut[13812] <= 16'd13529;
          lut[13813] <= 16'd13599;
          lut[13814] <= 16'd13668;
          lut[13815] <= 16'd13737;
          lut[13816] <= 16'd13805;
          lut[13817] <= 16'd13873;
          lut[13818] <= 16'd13940;
          lut[13819] <= 16'd14006;
          lut[13820] <= 16'd14072;
          lut[13821] <= 16'd14137;
          lut[13822] <= 16'd14201;
          lut[13823] <= 16'd14265;
          lut[13824] <= 0;
          lut[13825] <= 16'd152;
          lut[13826] <= 16'd303;
          lut[13827] <= 16'd455;
          lut[13828] <= 16'd607;
          lut[13829] <= 16'd758;
          lut[13830] <= 16'd909;
          lut[13831] <= 16'd1060;
          lut[13832] <= 16'd1211;
          lut[13833] <= 16'd1362;
          lut[13834] <= 16'd1513;
          lut[13835] <= 16'd1663;
          lut[13836] <= 16'd1813;
          lut[13837] <= 16'd1963;
          lut[13838] <= 16'd2112;
          lut[13839] <= 16'd2261;
          lut[13840] <= 16'd2410;
          lut[13841] <= 16'd2558;
          lut[13842] <= 16'd2706;
          lut[13843] <= 16'd2853;
          lut[13844] <= 16'd3000;
          lut[13845] <= 16'd3147;
          lut[13846] <= 16'd3292;
          lut[13847] <= 16'd3438;
          lut[13848] <= 16'd3583;
          lut[13849] <= 16'd3727;
          lut[13850] <= 16'd3871;
          lut[13851] <= 16'd4014;
          lut[13852] <= 16'd4156;
          lut[13853] <= 16'd4298;
          lut[13854] <= 16'd4439;
          lut[13855] <= 16'd4580;
          lut[13856] <= 16'd4720;
          lut[13857] <= 16'd4859;
          lut[13858] <= 16'd4997;
          lut[13859] <= 16'd5135;
          lut[13860] <= 16'd5272;
          lut[13861] <= 16'd5408;
          lut[13862] <= 16'd5543;
          lut[13863] <= 16'd5678;
          lut[13864] <= 16'd5811;
          lut[13865] <= 16'd5944;
          lut[13866] <= 16'd6077;
          lut[13867] <= 16'd6208;
          lut[13868] <= 16'd6339;
          lut[13869] <= 16'd6468;
          lut[13870] <= 16'd6597;
          lut[13871] <= 16'd6725;
          lut[13872] <= 16'd6852;
          lut[13873] <= 16'd6978;
          lut[13874] <= 16'd7104;
          lut[13875] <= 16'd7228;
          lut[13876] <= 16'd7352;
          lut[13877] <= 16'd7475;
          lut[13878] <= 16'd7596;
          lut[13879] <= 16'd7717;
          lut[13880] <= 16'd7837;
          lut[13881] <= 16'd7956;
          lut[13882] <= 16'd8075;
          lut[13883] <= 16'd8192;
          lut[13884] <= 16'd8308;
          lut[13885] <= 16'd8424;
          lut[13886] <= 16'd8538;
          lut[13887] <= 16'd8652;
          lut[13888] <= 16'd8765;
          lut[13889] <= 16'd8877;
          lut[13890] <= 16'd8987;
          lut[13891] <= 16'd9097;
          lut[13892] <= 16'd9207;
          lut[13893] <= 16'd9315;
          lut[13894] <= 16'd9422;
          lut[13895] <= 16'd9528;
          lut[13896] <= 16'd9634;
          lut[13897] <= 16'd9738;
          lut[13898] <= 16'd9842;
          lut[13899] <= 16'd9945;
          lut[13900] <= 16'd10047;
          lut[13901] <= 16'd10148;
          lut[13902] <= 16'd10248;
          lut[13903] <= 16'd10347;
          lut[13904] <= 16'd10446;
          lut[13905] <= 16'd10543;
          lut[13906] <= 16'd10640;
          lut[13907] <= 16'd10736;
          lut[13908] <= 16'd10831;
          lut[13909] <= 16'd10925;
          lut[13910] <= 16'd11018;
          lut[13911] <= 16'd11110;
          lut[13912] <= 16'd11202;
          lut[13913] <= 16'd11293;
          lut[13914] <= 16'd11383;
          lut[13915] <= 16'd11472;
          lut[13916] <= 16'd11560;
          lut[13917] <= 16'd11648;
          lut[13918] <= 16'd11734;
          lut[13919] <= 16'd11820;
          lut[13920] <= 16'd11905;
          lut[13921] <= 16'd11990;
          lut[13922] <= 16'd12073;
          lut[13923] <= 16'd12156;
          lut[13924] <= 16'd12238;
          lut[13925] <= 16'd12319;
          lut[13926] <= 16'd12400;
          lut[13927] <= 16'd12480;
          lut[13928] <= 16'd12559;
          lut[13929] <= 16'd12637;
          lut[13930] <= 16'd12715;
          lut[13931] <= 16'd12792;
          lut[13932] <= 16'd12868;
          lut[13933] <= 16'd12943;
          lut[13934] <= 16'd13018;
          lut[13935] <= 16'd13092;
          lut[13936] <= 16'd13166;
          lut[13937] <= 16'd13239;
          lut[13938] <= 16'd13311;
          lut[13939] <= 16'd13382;
          lut[13940] <= 16'd13453;
          lut[13941] <= 16'd13523;
          lut[13942] <= 16'd13592;
          lut[13943] <= 16'd13661;
          lut[13944] <= 16'd13729;
          lut[13945] <= 16'd13797;
          lut[13946] <= 16'd13864;
          lut[13947] <= 16'd13930;
          lut[13948] <= 16'd13996;
          lut[13949] <= 16'd14061;
          lut[13950] <= 16'd14126;
          lut[13951] <= 16'd14190;
          lut[13952] <= 0;
          lut[13953] <= 16'd150;
          lut[13954] <= 16'd301;
          lut[13955] <= 16'd451;
          lut[13956] <= 16'd601;
          lut[13957] <= 16'd751;
          lut[13958] <= 16'd901;
          lut[13959] <= 16'd1051;
          lut[13960] <= 16'd1200;
          lut[13961] <= 16'd1350;
          lut[13962] <= 16'd1499;
          lut[13963] <= 16'd1648;
          lut[13964] <= 16'd1797;
          lut[13965] <= 16'd1945;
          lut[13966] <= 16'd2093;
          lut[13967] <= 16'd2241;
          lut[13968] <= 16'd2388;
          lut[13969] <= 16'd2535;
          lut[13970] <= 16'd2681;
          lut[13971] <= 16'd2828;
          lut[13972] <= 16'd2973;
          lut[13973] <= 16'd3118;
          lut[13974] <= 16'd3263;
          lut[13975] <= 16'd3407;
          lut[13976] <= 16'd3551;
          lut[13977] <= 16'd3694;
          lut[13978] <= 16'd3836;
          lut[13979] <= 16'd3978;
          lut[13980] <= 16'd4120;
          lut[13981] <= 16'd4260;
          lut[13982] <= 16'd4400;
          lut[13983] <= 16'd4540;
          lut[13984] <= 16'd4679;
          lut[13985] <= 16'd4817;
          lut[13986] <= 16'd4954;
          lut[13987] <= 16'd5091;
          lut[13988] <= 16'd5226;
          lut[13989] <= 16'd5362;
          lut[13990] <= 16'd5496;
          lut[13991] <= 16'd5630;
          lut[13992] <= 16'd5762;
          lut[13993] <= 16'd5895;
          lut[13994] <= 16'd6026;
          lut[13995] <= 16'd6156;
          lut[13996] <= 16'd6286;
          lut[13997] <= 16'd6415;
          lut[13998] <= 16'd6543;
          lut[13999] <= 16'd6670;
          lut[14000] <= 16'd6796;
          lut[14001] <= 16'd6922;
          lut[14002] <= 16'd7046;
          lut[14003] <= 16'd7170;
          lut[14004] <= 16'd7293;
          lut[14005] <= 16'd7415;
          lut[14006] <= 16'd7536;
          lut[14007] <= 16'd7656;
          lut[14008] <= 16'd7776;
          lut[14009] <= 16'd7894;
          lut[14010] <= 16'd8012;
          lut[14011] <= 16'd8129;
          lut[14012] <= 16'd8244;
          lut[14013] <= 16'd8359;
          lut[14014] <= 16'd8473;
          lut[14015] <= 16'd8586;
          lut[14016] <= 16'd8699;
          lut[14017] <= 16'd8810;
          lut[14018] <= 16'd8920;
          lut[14019] <= 16'd9030;
          lut[14020] <= 16'd9139;
          lut[14021] <= 16'd9246;
          lut[14022] <= 16'd9353;
          lut[14023] <= 16'd9459;
          lut[14024] <= 16'd9564;
          lut[14025] <= 16'd9668;
          lut[14026] <= 16'd9772;
          lut[14027] <= 16'd9874;
          lut[14028] <= 16'd9976;
          lut[14029] <= 16'd10077;
          lut[14030] <= 16'd10176;
          lut[14031] <= 16'd10275;
          lut[14032] <= 16'd10373;
          lut[14033] <= 16'd10471;
          lut[14034] <= 16'd10567;
          lut[14035] <= 16'd10663;
          lut[14036] <= 16'd10757;
          lut[14037] <= 16'd10851;
          lut[14038] <= 16'd10944;
          lut[14039] <= 16'd11037;
          lut[14040] <= 16'd11128;
          lut[14041] <= 16'd11219;
          lut[14042] <= 16'd11308;
          lut[14043] <= 16'd11397;
          lut[14044] <= 16'd11486;
          lut[14045] <= 16'd11573;
          lut[14046] <= 16'd11660;
          lut[14047] <= 16'd11745;
          lut[14048] <= 16'd11830;
          lut[14049] <= 16'd11915;
          lut[14050] <= 16'd11998;
          lut[14051] <= 16'd12081;
          lut[14052] <= 16'd12163;
          lut[14053] <= 16'd12244;
          lut[14054] <= 16'd12325;
          lut[14055] <= 16'd12404;
          lut[14056] <= 16'd12483;
          lut[14057] <= 16'd12562;
          lut[14058] <= 16'd12639;
          lut[14059] <= 16'd12716;
          lut[14060] <= 16'd12792;
          lut[14061] <= 16'd12868;
          lut[14062] <= 16'd12943;
          lut[14063] <= 16'd13017;
          lut[14064] <= 16'd13090;
          lut[14065] <= 16'd13163;
          lut[14066] <= 16'd13235;
          lut[14067] <= 16'd13307;
          lut[14068] <= 16'd13378;
          lut[14069] <= 16'd13448;
          lut[14070] <= 16'd13517;
          lut[14071] <= 16'd13586;
          lut[14072] <= 16'd13654;
          lut[14073] <= 16'd13722;
          lut[14074] <= 16'd13789;
          lut[14075] <= 16'd13855;
          lut[14076] <= 16'd13921;
          lut[14077] <= 16'd13986;
          lut[14078] <= 16'd14051;
          lut[14079] <= 16'd14115;
          lut[14080] <= 0;
          lut[14081] <= 16'd149;
          lut[14082] <= 16'd298;
          lut[14083] <= 16'd447;
          lut[14084] <= 16'd596;
          lut[14085] <= 16'd744;
          lut[14086] <= 16'd893;
          lut[14087] <= 16'd1041;
          lut[14088] <= 16'd1189;
          lut[14089] <= 16'd1338;
          lut[14090] <= 16'd1485;
          lut[14091] <= 16'd1633;
          lut[14092] <= 16'd1780;
          lut[14093] <= 16'd1927;
          lut[14094] <= 16'd2074;
          lut[14095] <= 16'd2220;
          lut[14096] <= 16'd2367;
          lut[14097] <= 16'd2512;
          lut[14098] <= 16'd2657;
          lut[14099] <= 16'd2802;
          lut[14100] <= 16'd2947;
          lut[14101] <= 16'd3091;
          lut[14102] <= 16'd3234;
          lut[14103] <= 16'd3377;
          lut[14104] <= 16'd3520;
          lut[14105] <= 16'd3661;
          lut[14106] <= 16'd3803;
          lut[14107] <= 16'd3944;
          lut[14108] <= 16'd4084;
          lut[14109] <= 16'd4223;
          lut[14110] <= 16'd4362;
          lut[14111] <= 16'd4501;
          lut[14112] <= 16'd4638;
          lut[14113] <= 16'd4775;
          lut[14114] <= 16'd4912;
          lut[14115] <= 16'd5047;
          lut[14116] <= 16'd5182;
          lut[14117] <= 16'd5316;
          lut[14118] <= 16'd5450;
          lut[14119] <= 16'd5582;
          lut[14120] <= 16'd5714;
          lut[14121] <= 16'd5845;
          lut[14122] <= 16'd5976;
          lut[14123] <= 16'd6105;
          lut[14124] <= 16'd6234;
          lut[14125] <= 16'd6362;
          lut[14126] <= 16'd6489;
          lut[14127] <= 16'd6616;
          lut[14128] <= 16'd6741;
          lut[14129] <= 16'd6866;
          lut[14130] <= 16'd6990;
          lut[14131] <= 16'd7113;
          lut[14132] <= 16'd7235;
          lut[14133] <= 16'd7356;
          lut[14134] <= 16'd7477;
          lut[14135] <= 16'd7596;
          lut[14136] <= 16'd7715;
          lut[14137] <= 16'd7833;
          lut[14138] <= 16'd7950;
          lut[14139] <= 16'd8066;
          lut[14140] <= 16'd8181;
          lut[14141] <= 16'd8296;
          lut[14142] <= 16'd8409;
          lut[14143] <= 16'd8522;
          lut[14144] <= 16'd8633;
          lut[14145] <= 16'd8744;
          lut[14146] <= 16'd8854;
          lut[14147] <= 16'd8963;
          lut[14148] <= 16'd9072;
          lut[14149] <= 16'd9179;
          lut[14150] <= 16'd9285;
          lut[14151] <= 16'd9391;
          lut[14152] <= 16'd9496;
          lut[14153] <= 16'd9599;
          lut[14154] <= 16'd9702;
          lut[14155] <= 16'd9804;
          lut[14156] <= 16'd9906;
          lut[14157] <= 16'd10006;
          lut[14158] <= 16'd10106;
          lut[14159] <= 16'd10204;
          lut[14160] <= 16'd10302;
          lut[14161] <= 16'd10399;
          lut[14162] <= 16'd10495;
          lut[14163] <= 16'd10591;
          lut[14164] <= 16'd10685;
          lut[14165] <= 16'd10779;
          lut[14166] <= 16'd10872;
          lut[14167] <= 16'd10964;
          lut[14168] <= 16'd11055;
          lut[14169] <= 16'd11145;
          lut[14170] <= 16'd11235;
          lut[14171] <= 16'd11324;
          lut[14172] <= 16'd11412;
          lut[14173] <= 16'd11499;
          lut[14174] <= 16'd11586;
          lut[14175] <= 16'd11671;
          lut[14176] <= 16'd11756;
          lut[14177] <= 16'd11840;
          lut[14178] <= 16'd11924;
          lut[14179] <= 16'd12006;
          lut[14180] <= 16'd12088;
          lut[14181] <= 16'd12170;
          lut[14182] <= 16'd12250;
          lut[14183] <= 16'd12330;
          lut[14184] <= 16'd12409;
          lut[14185] <= 16'd12487;
          lut[14186] <= 16'd12565;
          lut[14187] <= 16'd12641;
          lut[14188] <= 16'd12718;
          lut[14189] <= 16'd12793;
          lut[14190] <= 16'd12868;
          lut[14191] <= 16'd12942;
          lut[14192] <= 16'd13016;
          lut[14193] <= 16'd13088;
          lut[14194] <= 16'd13161;
          lut[14195] <= 16'd13232;
          lut[14196] <= 16'd13303;
          lut[14197] <= 16'd13373;
          lut[14198] <= 16'd13443;
          lut[14199] <= 16'd13512;
          lut[14200] <= 16'd13580;
          lut[14201] <= 16'd13648;
          lut[14202] <= 16'd13715;
          lut[14203] <= 16'd13781;
          lut[14204] <= 16'd13847;
          lut[14205] <= 16'd13912;
          lut[14206] <= 16'd13977;
          lut[14207] <= 16'd14041;
          lut[14208] <= 0;
          lut[14209] <= 16'd148;
          lut[14210] <= 16'd295;
          lut[14211] <= 16'd443;
          lut[14212] <= 16'd590;
          lut[14213] <= 16'd738;
          lut[14214] <= 16'd885;
          lut[14215] <= 16'd1032;
          lut[14216] <= 16'd1179;
          lut[14217] <= 16'd1326;
          lut[14218] <= 16'd1472;
          lut[14219] <= 16'd1618;
          lut[14220] <= 16'd1764;
          lut[14221] <= 16'd1910;
          lut[14222] <= 16'd2056;
          lut[14223] <= 16'd2201;
          lut[14224] <= 16'd2346;
          lut[14225] <= 16'd2490;
          lut[14226] <= 16'd2634;
          lut[14227] <= 16'd2778;
          lut[14228] <= 16'd2921;
          lut[14229] <= 16'd3063;
          lut[14230] <= 16'd3206;
          lut[14231] <= 16'd3348;
          lut[14232] <= 16'd3489;
          lut[14233] <= 16'd3630;
          lut[14234] <= 16'd3770;
          lut[14235] <= 16'd3909;
          lut[14236] <= 16'd4048;
          lut[14237] <= 16'd4187;
          lut[14238] <= 16'd4325;
          lut[14239] <= 16'd4462;
          lut[14240] <= 16'd4599;
          lut[14241] <= 16'd4735;
          lut[14242] <= 16'd4870;
          lut[14243] <= 16'd5004;
          lut[14244] <= 16'd5138;
          lut[14245] <= 16'd5272;
          lut[14246] <= 16'd5404;
          lut[14247] <= 16'd5536;
          lut[14248] <= 16'd5667;
          lut[14249] <= 16'd5797;
          lut[14250] <= 16'd5927;
          lut[14251] <= 16'd6055;
          lut[14252] <= 16'd6183;
          lut[14253] <= 16'd6310;
          lut[14254] <= 16'd6437;
          lut[14255] <= 16'd6562;
          lut[14256] <= 16'd6687;
          lut[14257] <= 16'd6811;
          lut[14258] <= 16'd6934;
          lut[14259] <= 16'd7056;
          lut[14260] <= 16'd7178;
          lut[14261] <= 16'd7299;
          lut[14262] <= 16'd7418;
          lut[14263] <= 16'd7537;
          lut[14264] <= 16'd7655;
          lut[14265] <= 16'd7773;
          lut[14266] <= 16'd7889;
          lut[14267] <= 16'd8004;
          lut[14268] <= 16'd8119;
          lut[14269] <= 16'd8233;
          lut[14270] <= 16'd8346;
          lut[14271] <= 16'd8458;
          lut[14272] <= 16'd8569;
          lut[14273] <= 16'd8679;
          lut[14274] <= 16'd8789;
          lut[14275] <= 16'd8898;
          lut[14276] <= 16'd9005;
          lut[14277] <= 16'd9112;
          lut[14278] <= 16'd9218;
          lut[14279] <= 16'd9323;
          lut[14280] <= 16'd9428;
          lut[14281] <= 16'd9531;
          lut[14282] <= 16'd9634;
          lut[14283] <= 16'd9736;
          lut[14284] <= 16'd9837;
          lut[14285] <= 16'd9937;
          lut[14286] <= 16'd10036;
          lut[14287] <= 16'd10134;
          lut[14288] <= 16'd10232;
          lut[14289] <= 16'd10328;
          lut[14290] <= 16'd10424;
          lut[14291] <= 16'd10519;
          lut[14292] <= 16'd10614;
          lut[14293] <= 16'd10707;
          lut[14294] <= 16'd10800;
          lut[14295] <= 16'd10892;
          lut[14296] <= 16'd10983;
          lut[14297] <= 16'd11073;
          lut[14298] <= 16'd11162;
          lut[14299] <= 16'd11251;
          lut[14300] <= 16'd11339;
          lut[14301] <= 16'd11426;
          lut[14302] <= 16'd11512;
          lut[14303] <= 16'd11598;
          lut[14304] <= 16'd11683;
          lut[14305] <= 16'd11767;
          lut[14306] <= 16'd11850;
          lut[14307] <= 16'd11933;
          lut[14308] <= 16'd12015;
          lut[14309] <= 16'd12096;
          lut[14310] <= 16'd12176;
          lut[14311] <= 16'd12256;
          lut[14312] <= 16'd12335;
          lut[14313] <= 16'd12413;
          lut[14314] <= 16'd12491;
          lut[14315] <= 16'd12567;
          lut[14316] <= 16'd12644;
          lut[14317] <= 16'd12719;
          lut[14318] <= 16'd12794;
          lut[14319] <= 16'd12868;
          lut[14320] <= 16'd12941;
          lut[14321] <= 16'd13014;
          lut[14322] <= 16'd13086;
          lut[14323] <= 16'd13158;
          lut[14324] <= 16'd13229;
          lut[14325] <= 16'd13299;
          lut[14326] <= 16'd13369;
          lut[14327] <= 16'd13438;
          lut[14328] <= 16'd13506;
          lut[14329] <= 16'd13574;
          lut[14330] <= 16'd13641;
          lut[14331] <= 16'd13707;
          lut[14332] <= 16'd13773;
          lut[14333] <= 16'd13839;
          lut[14334] <= 16'd13904;
          lut[14335] <= 16'd13968;
          lut[14336] <= 0;
          lut[14337] <= 16'd146;
          lut[14338] <= 16'd293;
          lut[14339] <= 16'd439;
          lut[14340] <= 16'd585;
          lut[14341] <= 16'd731;
          lut[14342] <= 16'd877;
          lut[14343] <= 16'd1023;
          lut[14344] <= 16'd1168;
          lut[14345] <= 16'd1314;
          lut[14346] <= 16'd1459;
          lut[14347] <= 16'd1604;
          lut[14348] <= 16'd1749;
          lut[14349] <= 16'd1893;
          lut[14350] <= 16'd2037;
          lut[14351] <= 16'd2181;
          lut[14352] <= 16'd2325;
          lut[14353] <= 16'd2468;
          lut[14354] <= 16'd2611;
          lut[14355] <= 16'd2753;
          lut[14356] <= 16'd2895;
          lut[14357] <= 16'd3037;
          lut[14358] <= 16'd3178;
          lut[14359] <= 16'd3318;
          lut[14360] <= 16'd3459;
          lut[14361] <= 16'd3598;
          lut[14362] <= 16'd3737;
          lut[14363] <= 16'd3876;
          lut[14364] <= 16'd4014;
          lut[14365] <= 16'd4151;
          lut[14366] <= 16'd4288;
          lut[14367] <= 16'd4424;
          lut[14368] <= 16'd4560;
          lut[14369] <= 16'd4695;
          lut[14370] <= 16'd4829;
          lut[14371] <= 16'd4962;
          lut[14372] <= 16'd5095;
          lut[14373] <= 16'd5228;
          lut[14374] <= 16'd5359;
          lut[14375] <= 16'd5490;
          lut[14376] <= 16'd5620;
          lut[14377] <= 16'd5749;
          lut[14378] <= 16'd5878;
          lut[14379] <= 16'd6006;
          lut[14380] <= 16'd6133;
          lut[14381] <= 16'd6259;
          lut[14382] <= 16'd6385;
          lut[14383] <= 16'd6510;
          lut[14384] <= 16'd6634;
          lut[14385] <= 16'd6757;
          lut[14386] <= 16'd6879;
          lut[14387] <= 16'd7001;
          lut[14388] <= 16'd7122;
          lut[14389] <= 16'd7242;
          lut[14390] <= 16'd7361;
          lut[14391] <= 16'd7479;
          lut[14392] <= 16'd7596;
          lut[14393] <= 16'd7713;
          lut[14394] <= 16'd7829;
          lut[14395] <= 16'd7944;
          lut[14396] <= 16'd8058;
          lut[14397] <= 16'd8171;
          lut[14398] <= 16'd8283;
          lut[14399] <= 16'd8395;
          lut[14400] <= 16'd8506;
          lut[14401] <= 16'd8616;
          lut[14402] <= 16'd8725;
          lut[14403] <= 16'd8833;
          lut[14404] <= 16'd8940;
          lut[14405] <= 16'd9046;
          lut[14406] <= 16'd9152;
          lut[14407] <= 16'd9257;
          lut[14408] <= 16'd9361;
          lut[14409] <= 16'd9464;
          lut[14410] <= 16'd9566;
          lut[14411] <= 16'd9668;
          lut[14412] <= 16'd9768;
          lut[14413] <= 16'd9868;
          lut[14414] <= 16'd9967;
          lut[14415] <= 16'd10065;
          lut[14416] <= 16'd10162;
          lut[14417] <= 16'd10259;
          lut[14418] <= 16'd10354;
          lut[14419] <= 16'd10449;
          lut[14420] <= 16'd10543;
          lut[14421] <= 16'd10636;
          lut[14422] <= 16'd10729;
          lut[14423] <= 16'd10820;
          lut[14424] <= 16'd10911;
          lut[14425] <= 16'd11001;
          lut[14426] <= 16'd11091;
          lut[14427] <= 16'd11179;
          lut[14428] <= 16'd11267;
          lut[14429] <= 16'd11354;
          lut[14430] <= 16'd11440;
          lut[14431] <= 16'd11525;
          lut[14432] <= 16'd11610;
          lut[14433] <= 16'd11694;
          lut[14434] <= 16'd11777;
          lut[14435] <= 16'd11860;
          lut[14436] <= 16'd11942;
          lut[14437] <= 16'd12023;
          lut[14438] <= 16'd12103;
          lut[14439] <= 16'd12183;
          lut[14440] <= 16'd12261;
          lut[14441] <= 16'd12340;
          lut[14442] <= 16'd12417;
          lut[14443] <= 16'd12494;
          lut[14444] <= 16'd12570;
          lut[14445] <= 16'd12646;
          lut[14446] <= 16'd12720;
          lut[14447] <= 16'd12794;
          lut[14448] <= 16'd12868;
          lut[14449] <= 16'd12941;
          lut[14450] <= 16'd13013;
          lut[14451] <= 16'd13084;
          lut[14452] <= 16'd13155;
          lut[14453] <= 16'd13226;
          lut[14454] <= 16'd13295;
          lut[14455] <= 16'd13364;
          lut[14456] <= 16'd13433;
          lut[14457] <= 16'd13501;
          lut[14458] <= 16'd13568;
          lut[14459] <= 16'd13634;
          lut[14460] <= 16'd13700;
          lut[14461] <= 16'd13766;
          lut[14462] <= 16'd13831;
          lut[14463] <= 16'd13895;
          lut[14464] <= 0;
          lut[14465] <= 16'd145;
          lut[14466] <= 16'd290;
          lut[14467] <= 16'd435;
          lut[14468] <= 16'd580;
          lut[14469] <= 16'd724;
          lut[14470] <= 16'd869;
          lut[14471] <= 16'd1014;
          lut[14472] <= 16'd1158;
          lut[14473] <= 16'd1302;
          lut[14474] <= 16'd1446;
          lut[14475] <= 16'd1590;
          lut[14476] <= 16'd1733;
          lut[14477] <= 16'd1877;
          lut[14478] <= 16'd2020;
          lut[14479] <= 16'd2162;
          lut[14480] <= 16'd2305;
          lut[14481] <= 16'd2447;
          lut[14482] <= 16'd2588;
          lut[14483] <= 16'd2729;
          lut[14484] <= 16'd2870;
          lut[14485] <= 16'd3010;
          lut[14486] <= 16'd3150;
          lut[14487] <= 16'd3290;
          lut[14488] <= 16'd3429;
          lut[14489] <= 16'd3567;
          lut[14490] <= 16'd3705;
          lut[14491] <= 16'd3843;
          lut[14492] <= 16'd3980;
          lut[14493] <= 16'd4116;
          lut[14494] <= 16'd4252;
          lut[14495] <= 16'd4387;
          lut[14496] <= 16'd4521;
          lut[14497] <= 16'd4655;
          lut[14498] <= 16'd4789;
          lut[14499] <= 16'd4921;
          lut[14500] <= 16'd5053;
          lut[14501] <= 16'd5184;
          lut[14502] <= 16'd5315;
          lut[14503] <= 16'd5445;
          lut[14504] <= 16'd5574;
          lut[14505] <= 16'd5703;
          lut[14506] <= 16'd5830;
          lut[14507] <= 16'd5957;
          lut[14508] <= 16'd6084;
          lut[14509] <= 16'd6209;
          lut[14510] <= 16'd6334;
          lut[14511] <= 16'd6458;
          lut[14512] <= 16'd6581;
          lut[14513] <= 16'd6704;
          lut[14514] <= 16'd6825;
          lut[14515] <= 16'd6946;
          lut[14516] <= 16'd7066;
          lut[14517] <= 16'd7185;
          lut[14518] <= 16'd7304;
          lut[14519] <= 16'd7421;
          lut[14520] <= 16'd7538;
          lut[14521] <= 16'd7654;
          lut[14522] <= 16'd7769;
          lut[14523] <= 16'd7884;
          lut[14524] <= 16'd7997;
          lut[14525] <= 16'd8110;
          lut[14526] <= 16'd8222;
          lut[14527] <= 16'd8333;
          lut[14528] <= 16'd8443;
          lut[14529] <= 16'd8552;
          lut[14530] <= 16'd8661;
          lut[14531] <= 16'd8769;
          lut[14532] <= 16'd8876;
          lut[14533] <= 16'd8982;
          lut[14534] <= 16'd9087;
          lut[14535] <= 16'd9191;
          lut[14536] <= 16'd9295;
          lut[14537] <= 16'd9397;
          lut[14538] <= 16'd9499;
          lut[14539] <= 16'd9600;
          lut[14540] <= 16'd9701;
          lut[14541] <= 16'd9800;
          lut[14542] <= 16'd9899;
          lut[14543] <= 16'd9996;
          lut[14544] <= 16'd10093;
          lut[14545] <= 16'd10190;
          lut[14546] <= 16'd10285;
          lut[14547] <= 16'd10380;
          lut[14548] <= 16'd10473;
          lut[14549] <= 16'd10566;
          lut[14550] <= 16'd10659;
          lut[14551] <= 16'd10750;
          lut[14552] <= 16'd10841;
          lut[14553] <= 16'd10930;
          lut[14554] <= 16'd11020;
          lut[14555] <= 16'd11108;
          lut[14556] <= 16'd11195;
          lut[14557] <= 16'd11282;
          lut[14558] <= 16'd11368;
          lut[14559] <= 16'd11454;
          lut[14560] <= 16'd11538;
          lut[14561] <= 16'd11622;
          lut[14562] <= 16'd11705;
          lut[14563] <= 16'd11788;
          lut[14564] <= 16'd11869;
          lut[14565] <= 16'd11950;
          lut[14566] <= 16'd12030;
          lut[14567] <= 16'd12110;
          lut[14568] <= 16'd12189;
          lut[14569] <= 16'd12267;
          lut[14570] <= 16'd12344;
          lut[14571] <= 16'd12421;
          lut[14572] <= 16'd12497;
          lut[14573] <= 16'd12573;
          lut[14574] <= 16'd12648;
          lut[14575] <= 16'd12722;
          lut[14576] <= 16'd12795;
          lut[14577] <= 16'd12868;
          lut[14578] <= 16'd12940;
          lut[14579] <= 16'd13012;
          lut[14580] <= 16'd13083;
          lut[14581] <= 16'd13153;
          lut[14582] <= 16'd13223;
          lut[14583] <= 16'd13292;
          lut[14584] <= 16'd13360;
          lut[14585] <= 16'd13428;
          lut[14586] <= 16'd13495;
          lut[14587] <= 16'd13562;
          lut[14588] <= 16'd13628;
          lut[14589] <= 16'd13693;
          lut[14590] <= 16'd13758;
          lut[14591] <= 16'd13823;
          lut[14592] <= 0;
          lut[14593] <= 16'd144;
          lut[14594] <= 16'd287;
          lut[14595] <= 16'd431;
          lut[14596] <= 16'd575;
          lut[14597] <= 16'd718;
          lut[14598] <= 16'd862;
          lut[14599] <= 16'd1005;
          lut[14600] <= 16'd1148;
          lut[14601] <= 16'd1291;
          lut[14602] <= 16'd1434;
          lut[14603] <= 16'd1576;
          lut[14604] <= 16'd1718;
          lut[14605] <= 16'd1860;
          lut[14606] <= 16'd2002;
          lut[14607] <= 16'd2143;
          lut[14608] <= 16'd2285;
          lut[14609] <= 16'd2425;
          lut[14610] <= 16'd2566;
          lut[14611] <= 16'd2706;
          lut[14612] <= 16'd2845;
          lut[14613] <= 16'd2985;
          lut[14614] <= 16'd3123;
          lut[14615] <= 16'd3262;
          lut[14616] <= 16'd3400;
          lut[14617] <= 16'd3537;
          lut[14618] <= 16'd3674;
          lut[14619] <= 16'd3810;
          lut[14620] <= 16'd3946;
          lut[14621] <= 16'd4081;
          lut[14622] <= 16'd4216;
          lut[14623] <= 16'd4350;
          lut[14624] <= 16'd4484;
          lut[14625] <= 16'd4617;
          lut[14626] <= 16'd4749;
          lut[14627] <= 16'd4881;
          lut[14628] <= 16'd5012;
          lut[14629] <= 16'd5142;
          lut[14630] <= 16'd5272;
          lut[14631] <= 16'd5401;
          lut[14632] <= 16'd5529;
          lut[14633] <= 16'd5656;
          lut[14634] <= 16'd5783;
          lut[14635] <= 16'd5910;
          lut[14636] <= 16'd6035;
          lut[14637] <= 16'd6160;
          lut[14638] <= 16'd6284;
          lut[14639] <= 16'd6407;
          lut[14640] <= 16'd6529;
          lut[14641] <= 16'd6651;
          lut[14642] <= 16'd6772;
          lut[14643] <= 16'd6892;
          lut[14644] <= 16'd7012;
          lut[14645] <= 16'd7130;
          lut[14646] <= 16'd7248;
          lut[14647] <= 16'd7365;
          lut[14648] <= 16'd7481;
          lut[14649] <= 16'd7596;
          lut[14650] <= 16'd7711;
          lut[14651] <= 16'd7825;
          lut[14652] <= 16'd7938;
          lut[14653] <= 16'd8050;
          lut[14654] <= 16'd8161;
          lut[14655] <= 16'd8272;
          lut[14656] <= 16'd8381;
          lut[14657] <= 16'd8490;
          lut[14658] <= 16'd8598;
          lut[14659] <= 16'd8705;
          lut[14660] <= 16'd8812;
          lut[14661] <= 16'd8917;
          lut[14662] <= 16'd9022;
          lut[14663] <= 16'd9126;
          lut[14664] <= 16'd9229;
          lut[14665] <= 16'd9332;
          lut[14666] <= 16'd9433;
          lut[14667] <= 16'd9534;
          lut[14668] <= 16'd9634;
          lut[14669] <= 16'd9733;
          lut[14670] <= 16'd9831;
          lut[14671] <= 16'd9929;
          lut[14672] <= 16'd10025;
          lut[14673] <= 16'd10121;
          lut[14674] <= 16'd10216;
          lut[14675] <= 16'd10311;
          lut[14676] <= 16'd10404;
          lut[14677] <= 16'd10497;
          lut[14678] <= 16'd10589;
          lut[14679] <= 16'd10680;
          lut[14680] <= 16'd10771;
          lut[14681] <= 16'd10860;
          lut[14682] <= 16'd10949;
          lut[14683] <= 16'd11037;
          lut[14684] <= 16'd11125;
          lut[14685] <= 16'd11211;
          lut[14686] <= 16'd11297;
          lut[14687] <= 16'd11383;
          lut[14688] <= 16'd11467;
          lut[14689] <= 16'd11551;
          lut[14690] <= 16'd11634;
          lut[14691] <= 16'd11716;
          lut[14692] <= 16'd11798;
          lut[14693] <= 16'd11879;
          lut[14694] <= 16'd11959;
          lut[14695] <= 16'd12038;
          lut[14696] <= 16'd12117;
          lut[14697] <= 16'd12195;
          lut[14698] <= 16'd12272;
          lut[14699] <= 16'd12349;
          lut[14700] <= 16'd12425;
          lut[14701] <= 16'd12501;
          lut[14702] <= 16'd12575;
          lut[14703] <= 16'd12650;
          lut[14704] <= 16'd12723;
          lut[14705] <= 16'd12796;
          lut[14706] <= 16'd12868;
          lut[14707] <= 16'd12940;
          lut[14708] <= 16'd13010;
          lut[14709] <= 16'd13081;
          lut[14710] <= 16'd13150;
          lut[14711] <= 16'd13219;
          lut[14712] <= 16'd13288;
          lut[14713] <= 16'd13356;
          lut[14714] <= 16'd13423;
          lut[14715] <= 16'd13490;
          lut[14716] <= 16'd13556;
          lut[14717] <= 16'd13622;
          lut[14718] <= 16'd13686;
          lut[14719] <= 16'd13751;
          lut[14720] <= 0;
          lut[14721] <= 16'd142;
          lut[14722] <= 16'd285;
          lut[14723] <= 16'd427;
          lut[14724] <= 16'd570;
          lut[14725] <= 16'd712;
          lut[14726] <= 16'd854;
          lut[14727] <= 16'd996;
          lut[14728] <= 16'd1138;
          lut[14729] <= 16'd1280;
          lut[14730] <= 16'd1421;
          lut[14731] <= 16'd1562;
          lut[14732] <= 16'd1703;
          lut[14733] <= 16'd1844;
          lut[14734] <= 16'd1985;
          lut[14735] <= 16'd2125;
          lut[14736] <= 16'd2265;
          lut[14737] <= 16'd2405;
          lut[14738] <= 16'd2544;
          lut[14739] <= 16'd2683;
          lut[14740] <= 16'd2821;
          lut[14741] <= 16'd2959;
          lut[14742] <= 16'd3097;
          lut[14743] <= 16'd3234;
          lut[14744] <= 16'd3371;
          lut[14745] <= 16'd3507;
          lut[14746] <= 16'd3643;
          lut[14747] <= 16'd3778;
          lut[14748] <= 16'd3913;
          lut[14749] <= 16'd4047;
          lut[14750] <= 16'd4181;
          lut[14751] <= 16'd4314;
          lut[14752] <= 16'd4447;
          lut[14753] <= 16'd4578;
          lut[14754] <= 16'd4710;
          lut[14755] <= 16'd4841;
          lut[14756] <= 16'd4971;
          lut[14757] <= 16'd5100;
          lut[14758] <= 16'd5229;
          lut[14759] <= 16'd5357;
          lut[14760] <= 16'd5484;
          lut[14761] <= 16'd5611;
          lut[14762] <= 16'd5737;
          lut[14763] <= 16'd5862;
          lut[14764] <= 16'd5987;
          lut[14765] <= 16'd6111;
          lut[14766] <= 16'd6234;
          lut[14767] <= 16'd6357;
          lut[14768] <= 16'd6478;
          lut[14769] <= 16'd6599;
          lut[14770] <= 16'd6720;
          lut[14771] <= 16'd6839;
          lut[14772] <= 16'd6958;
          lut[14773] <= 16'd7076;
          lut[14774] <= 16'd7193;
          lut[14775] <= 16'd7309;
          lut[14776] <= 16'd7425;
          lut[14777] <= 16'd7539;
          lut[14778] <= 16'd7653;
          lut[14779] <= 16'd7766;
          lut[14780] <= 16'd7879;
          lut[14781] <= 16'd7990;
          lut[14782] <= 16'd8101;
          lut[14783] <= 16'd8211;
          lut[14784] <= 16'd8320;
          lut[14785] <= 16'd8429;
          lut[14786] <= 16'd8536;
          lut[14787] <= 16'd8643;
          lut[14788] <= 16'd8749;
          lut[14789] <= 16'd8854;
          lut[14790] <= 16'd8959;
          lut[14791] <= 16'd9062;
          lut[14792] <= 16'd9165;
          lut[14793] <= 16'd9267;
          lut[14794] <= 16'd9368;
          lut[14795] <= 16'd9468;
          lut[14796] <= 16'd9568;
          lut[14797] <= 16'd9667;
          lut[14798] <= 16'd9765;
          lut[14799] <= 16'd9862;
          lut[14800] <= 16'd9958;
          lut[14801] <= 16'd10054;
          lut[14802] <= 16'd10149;
          lut[14803] <= 16'd10243;
          lut[14804] <= 16'd10336;
          lut[14805] <= 16'd10429;
          lut[14806] <= 16'd10520;
          lut[14807] <= 16'd10611;
          lut[14808] <= 16'd10702;
          lut[14809] <= 16'd10791;
          lut[14810] <= 16'd10880;
          lut[14811] <= 16'd10968;
          lut[14812] <= 16'd11055;
          lut[14813] <= 16'd11141;
          lut[14814] <= 16'd11227;
          lut[14815] <= 16'd11312;
          lut[14816] <= 16'd11397;
          lut[14817] <= 16'd11480;
          lut[14818] <= 16'd11563;
          lut[14819] <= 16'd11645;
          lut[14820] <= 16'd11727;
          lut[14821] <= 16'd11808;
          lut[14822] <= 16'd11888;
          lut[14823] <= 16'd11967;
          lut[14824] <= 16'd12046;
          lut[14825] <= 16'd12124;
          lut[14826] <= 16'd12201;
          lut[14827] <= 16'd12278;
          lut[14828] <= 16'd12354;
          lut[14829] <= 16'd12429;
          lut[14830] <= 16'd12504;
          lut[14831] <= 16'd12578;
          lut[14832] <= 16'd12651;
          lut[14833] <= 16'd12724;
          lut[14834] <= 16'd12796;
          lut[14835] <= 16'd12868;
          lut[14836] <= 16'd12939;
          lut[14837] <= 16'd13009;
          lut[14838] <= 16'd13079;
          lut[14839] <= 16'd13148;
          lut[14840] <= 16'd13217;
          lut[14841] <= 16'd13284;
          lut[14842] <= 16'd13352;
          lut[14843] <= 16'd13418;
          lut[14844] <= 16'd13485;
          lut[14845] <= 16'd13550;
          lut[14846] <= 16'd13615;
          lut[14847] <= 16'd13680;
          lut[14848] <= 0;
          lut[14849] <= 16'd141;
          lut[14850] <= 16'd282;
          lut[14851] <= 16'd424;
          lut[14852] <= 16'd565;
          lut[14853] <= 16'd706;
          lut[14854] <= 16'd847;
          lut[14855] <= 16'd987;
          lut[14856] <= 16'd1128;
          lut[14857] <= 16'd1269;
          lut[14858] <= 16'd1409;
          lut[14859] <= 16'd1549;
          lut[14860] <= 16'd1689;
          lut[14861] <= 16'd1829;
          lut[14862] <= 16'd1968;
          lut[14863] <= 16'd2107;
          lut[14864] <= 16'd2246;
          lut[14865] <= 16'd2384;
          lut[14866] <= 16'd2522;
          lut[14867] <= 16'd2660;
          lut[14868] <= 16'd2797;
          lut[14869] <= 16'd2934;
          lut[14870] <= 16'd3071;
          lut[14871] <= 16'd3207;
          lut[14872] <= 16'd3343;
          lut[14873] <= 16'd3478;
          lut[14874] <= 16'd3613;
          lut[14875] <= 16'd3747;
          lut[14876] <= 16'd3881;
          lut[14877] <= 16'd4014;
          lut[14878] <= 16'd4146;
          lut[14879] <= 16'd4278;
          lut[14880] <= 16'd4410;
          lut[14881] <= 16'd4541;
          lut[14882] <= 16'd4671;
          lut[14883] <= 16'd4801;
          lut[14884] <= 16'd4930;
          lut[14885] <= 16'd5059;
          lut[14886] <= 16'd5187;
          lut[14887] <= 16'd5314;
          lut[14888] <= 16'd5440;
          lut[14889] <= 16'd5566;
          lut[14890] <= 16'd5692;
          lut[14891] <= 16'd5816;
          lut[14892] <= 16'd5940;
          lut[14893] <= 16'd6063;
          lut[14894] <= 16'd6185;
          lut[14895] <= 16'd6307;
          lut[14896] <= 16'd6428;
          lut[14897] <= 16'd6548;
          lut[14898] <= 16'd6668;
          lut[14899] <= 16'd6787;
          lut[14900] <= 16'd6905;
          lut[14901] <= 16'd7022;
          lut[14902] <= 16'd7138;
          lut[14903] <= 16'd7254;
          lut[14904] <= 16'd7369;
          lut[14905] <= 16'd7483;
          lut[14906] <= 16'd7596;
          lut[14907] <= 16'd7709;
          lut[14908] <= 16'd7821;
          lut[14909] <= 16'd7932;
          lut[14910] <= 16'd8042;
          lut[14911] <= 16'd8152;
          lut[14912] <= 16'd8260;
          lut[14913] <= 16'd8368;
          lut[14914] <= 16'd8475;
          lut[14915] <= 16'd8582;
          lut[14916] <= 16'd8687;
          lut[14917] <= 16'd8792;
          lut[14918] <= 16'd8896;
          lut[14919] <= 16'd8999;
          lut[14920] <= 16'd9101;
          lut[14921] <= 16'd9203;
          lut[14922] <= 16'd9304;
          lut[14923] <= 16'd9404;
          lut[14924] <= 16'd9503;
          lut[14925] <= 16'd9601;
          lut[14926] <= 16'd9699;
          lut[14927] <= 16'd9796;
          lut[14928] <= 16'd9892;
          lut[14929] <= 16'd9987;
          lut[14930] <= 16'd10082;
          lut[14931] <= 16'd10176;
          lut[14932] <= 16'd10269;
          lut[14933] <= 16'd10361;
          lut[14934] <= 16'd10452;
          lut[14935] <= 16'd10543;
          lut[14936] <= 16'd10633;
          lut[14937] <= 16'd10722;
          lut[14938] <= 16'd10811;
          lut[14939] <= 16'd10899;
          lut[14940] <= 16'd10986;
          lut[14941] <= 16'd11072;
          lut[14942] <= 16'd11158;
          lut[14943] <= 16'd11243;
          lut[14944] <= 16'd11327;
          lut[14945] <= 16'd11410;
          lut[14946] <= 16'd11493;
          lut[14947] <= 16'd11575;
          lut[14948] <= 16'd11657;
          lut[14949] <= 16'd11737;
          lut[14950] <= 16'd11817;
          lut[14951] <= 16'd11897;
          lut[14952] <= 16'd11975;
          lut[14953] <= 16'd12053;
          lut[14954] <= 16'd12130;
          lut[14955] <= 16'd12207;
          lut[14956] <= 16'd12283;
          lut[14957] <= 16'd12358;
          lut[14958] <= 16'd12433;
          lut[14959] <= 16'd12507;
          lut[14960] <= 16'd12581;
          lut[14961] <= 16'd12653;
          lut[14962] <= 16'd12725;
          lut[14963] <= 16'd12797;
          lut[14964] <= 16'd12868;
          lut[14965] <= 16'd12938;
          lut[14966] <= 16'd13008;
          lut[14967] <= 16'd13077;
          lut[14968] <= 16'd13146;
          lut[14969] <= 16'd13214;
          lut[14970] <= 16'd13281;
          lut[14971] <= 16'd13348;
          lut[14972] <= 16'd13414;
          lut[14973] <= 16'd13480;
          lut[14974] <= 16'd13545;
          lut[14975] <= 16'd13609;
          lut[14976] <= 0;
          lut[14977] <= 16'd140;
          lut[14978] <= 16'd280;
          lut[14979] <= 16'd420;
          lut[14980] <= 16'd560;
          lut[14981] <= 16'd700;
          lut[14982] <= 16'd839;
          lut[14983] <= 16'd979;
          lut[14984] <= 16'd1119;
          lut[14985] <= 16'd1258;
          lut[14986] <= 16'd1397;
          lut[14987] <= 16'd1536;
          lut[14988] <= 16'd1675;
          lut[14989] <= 16'd1813;
          lut[14990] <= 16'd1951;
          lut[14991] <= 16'd2089;
          lut[14992] <= 16'd2227;
          lut[14993] <= 16'd2364;
          lut[14994] <= 16'd2501;
          lut[14995] <= 16'd2638;
          lut[14996] <= 16'd2774;
          lut[14997] <= 16'd2910;
          lut[14998] <= 16'd3045;
          lut[14999] <= 16'd3180;
          lut[15000] <= 16'd3315;
          lut[15001] <= 16'd3449;
          lut[15002] <= 16'd3583;
          lut[15003] <= 16'd3716;
          lut[15004] <= 16'd3849;
          lut[15005] <= 16'd3981;
          lut[15006] <= 16'd4112;
          lut[15007] <= 16'd4244;
          lut[15008] <= 16'd4374;
          lut[15009] <= 16'd4504;
          lut[15010] <= 16'd4634;
          lut[15011] <= 16'd4762;
          lut[15012] <= 16'd4891;
          lut[15013] <= 16'd5018;
          lut[15014] <= 16'd5145;
          lut[15015] <= 16'd5272;
          lut[15016] <= 16'd5397;
          lut[15017] <= 16'd5522;
          lut[15018] <= 16'd5647;
          lut[15019] <= 16'd5770;
          lut[15020] <= 16'd5893;
          lut[15021] <= 16'd6016;
          lut[15022] <= 16'd6137;
          lut[15023] <= 16'd6258;
          lut[15024] <= 16'd6379;
          lut[15025] <= 16'd6498;
          lut[15026] <= 16'd6617;
          lut[15027] <= 16'd6735;
          lut[15028] <= 16'd6852;
          lut[15029] <= 16'd6969;
          lut[15030] <= 16'd7085;
          lut[15031] <= 16'd7200;
          lut[15032] <= 16'd7314;
          lut[15033] <= 16'd7428;
          lut[15034] <= 16'd7540;
          lut[15035] <= 16'd7652;
          lut[15036] <= 16'd7764;
          lut[15037] <= 16'd7874;
          lut[15038] <= 16'd7984;
          lut[15039] <= 16'd8093;
          lut[15040] <= 16'd8201;
          lut[15041] <= 16'd8308;
          lut[15042] <= 16'd8415;
          lut[15043] <= 16'd8521;
          lut[15044] <= 16'd8626;
          lut[15045] <= 16'd8730;
          lut[15046] <= 16'd8834;
          lut[15047] <= 16'd8936;
          lut[15048] <= 16'd9038;
          lut[15049] <= 16'd9139;
          lut[15050] <= 16'd9240;
          lut[15051] <= 16'd9340;
          lut[15052] <= 16'd9438;
          lut[15053] <= 16'd9537;
          lut[15054] <= 16'd9634;
          lut[15055] <= 16'd9730;
          lut[15056] <= 16'd9826;
          lut[15057] <= 16'd9921;
          lut[15058] <= 16'd10016;
          lut[15059] <= 16'd10109;
          lut[15060] <= 16'd10202;
          lut[15061] <= 16'd10294;
          lut[15062] <= 16'd10385;
          lut[15063] <= 16'd10476;
          lut[15064] <= 16'd10566;
          lut[15065] <= 16'd10655;
          lut[15066] <= 16'd10743;
          lut[15067] <= 16'd10831;
          lut[15068] <= 16'd10917;
          lut[15069] <= 16'd11004;
          lut[15070] <= 16'd11089;
          lut[15071] <= 16'd11174;
          lut[15072] <= 16'd11258;
          lut[15073] <= 16'd11341;
          lut[15074] <= 16'd11424;
          lut[15075] <= 16'd11506;
          lut[15076] <= 16'd11587;
          lut[15077] <= 16'd11668;
          lut[15078] <= 16'd11748;
          lut[15079] <= 16'd11827;
          lut[15080] <= 16'd11905;
          lut[15081] <= 16'd11983;
          lut[15082] <= 16'd12060;
          lut[15083] <= 16'd12137;
          lut[15084] <= 16'd12213;
          lut[15085] <= 16'd12288;
          lut[15086] <= 16'd12363;
          lut[15087] <= 16'd12437;
          lut[15088] <= 16'd12510;
          lut[15089] <= 16'd12583;
          lut[15090] <= 16'd12655;
          lut[15091] <= 16'd12727;
          lut[15092] <= 16'd12798;
          lut[15093] <= 16'd12868;
          lut[15094] <= 16'd12938;
          lut[15095] <= 16'd13007;
          lut[15096] <= 16'd13075;
          lut[15097] <= 16'd13143;
          lut[15098] <= 16'd13211;
          lut[15099] <= 16'd13277;
          lut[15100] <= 16'd13344;
          lut[15101] <= 16'd13409;
          lut[15102] <= 16'd13475;
          lut[15103] <= 16'd13539;
          lut[15104] <= 0;
          lut[15105] <= 16'd139;
          lut[15106] <= 16'd278;
          lut[15107] <= 16'd416;
          lut[15108] <= 16'd555;
          lut[15109] <= 16'd694;
          lut[15110] <= 16'd832;
          lut[15111] <= 16'd971;
          lut[15112] <= 16'd1109;
          lut[15113] <= 16'd1247;
          lut[15114] <= 16'd1385;
          lut[15115] <= 16'd1523;
          lut[15116] <= 16'd1660;
          lut[15117] <= 16'd1798;
          lut[15118] <= 16'd1935;
          lut[15119] <= 16'd2072;
          lut[15120] <= 16'd2208;
          lut[15121] <= 16'd2344;
          lut[15122] <= 16'd2480;
          lut[15123] <= 16'd2616;
          lut[15124] <= 16'd2751;
          lut[15125] <= 16'd2886;
          lut[15126] <= 16'd3020;
          lut[15127] <= 16'd3154;
          lut[15128] <= 16'd3287;
          lut[15129] <= 16'd3421;
          lut[15130] <= 16'd3553;
          lut[15131] <= 16'd3685;
          lut[15132] <= 16'd3817;
          lut[15133] <= 16'd3948;
          lut[15134] <= 16'd4079;
          lut[15135] <= 16'd4209;
          lut[15136] <= 16'd4339;
          lut[15137] <= 16'd4468;
          lut[15138] <= 16'd4596;
          lut[15139] <= 16'd4724;
          lut[15140] <= 16'd4852;
          lut[15141] <= 16'd4978;
          lut[15142] <= 16'd5104;
          lut[15143] <= 16'd5230;
          lut[15144] <= 16'd5355;
          lut[15145] <= 16'd5479;
          lut[15146] <= 16'd5603;
          lut[15147] <= 16'd5725;
          lut[15148] <= 16'd5848;
          lut[15149] <= 16'd5969;
          lut[15150] <= 16'd6090;
          lut[15151] <= 16'd6210;
          lut[15152] <= 16'd6330;
          lut[15153] <= 16'd6449;
          lut[15154] <= 16'd6567;
          lut[15155] <= 16'd6684;
          lut[15156] <= 16'd6801;
          lut[15157] <= 16'd6916;
          lut[15158] <= 16'd7032;
          lut[15159] <= 16'd7146;
          lut[15160] <= 16'd7260;
          lut[15161] <= 16'd7373;
          lut[15162] <= 16'd7485;
          lut[15163] <= 16'd7596;
          lut[15164] <= 16'd7707;
          lut[15165] <= 16'd7817;
          lut[15166] <= 16'd7926;
          lut[15167] <= 16'd8035;
          lut[15168] <= 16'd8142;
          lut[15169] <= 16'd8249;
          lut[15170] <= 16'd8355;
          lut[15171] <= 16'd8461;
          lut[15172] <= 16'd8565;
          lut[15173] <= 16'd8669;
          lut[15174] <= 16'd8772;
          lut[15175] <= 16'd8875;
          lut[15176] <= 16'd8976;
          lut[15177] <= 16'd9077;
          lut[15178] <= 16'd9177;
          lut[15179] <= 16'd9276;
          lut[15180] <= 16'd9375;
          lut[15181] <= 16'd9473;
          lut[15182] <= 16'd9570;
          lut[15183] <= 16'd9666;
          lut[15184] <= 16'd9761;
          lut[15185] <= 16'd9856;
          lut[15186] <= 16'd9950;
          lut[15187] <= 16'd10043;
          lut[15188] <= 16'd10136;
          lut[15189] <= 16'd10228;
          lut[15190] <= 16'd10319;
          lut[15191] <= 16'd10409;
          lut[15192] <= 16'd10499;
          lut[15193] <= 16'd10587;
          lut[15194] <= 16'd10676;
          lut[15195] <= 16'd10763;
          lut[15196] <= 16'd10850;
          lut[15197] <= 16'd10936;
          lut[15198] <= 16'd11021;
          lut[15199] <= 16'd11106;
          lut[15200] <= 16'd11190;
          lut[15201] <= 16'd11273;
          lut[15202] <= 16'd11355;
          lut[15203] <= 16'd11437;
          lut[15204] <= 16'd11518;
          lut[15205] <= 16'd11599;
          lut[15206] <= 16'd11678;
          lut[15207] <= 16'd11758;
          lut[15208] <= 16'd11836;
          lut[15209] <= 16'd11914;
          lut[15210] <= 16'd11991;
          lut[15211] <= 16'd12068;
          lut[15212] <= 16'd12143;
          lut[15213] <= 16'd12219;
          lut[15214] <= 16'd12293;
          lut[15215] <= 16'd12367;
          lut[15216] <= 16'd12441;
          lut[15217] <= 16'd12513;
          lut[15218] <= 16'd12586;
          lut[15219] <= 16'd12657;
          lut[15220] <= 16'd12728;
          lut[15221] <= 16'd12798;
          lut[15222] <= 16'd12868;
          lut[15223] <= 16'd12937;
          lut[15224] <= 16'd13006;
          lut[15225] <= 16'd13074;
          lut[15226] <= 16'd13141;
          lut[15227] <= 16'd13208;
          lut[15228] <= 16'd13274;
          lut[15229] <= 16'd13340;
          lut[15230] <= 16'd13405;
          lut[15231] <= 16'd13470;
          lut[15232] <= 0;
          lut[15233] <= 16'd138;
          lut[15234] <= 16'd275;
          lut[15235] <= 16'd413;
          lut[15236] <= 16'd551;
          lut[15237] <= 16'd688;
          lut[15238] <= 16'd825;
          lut[15239] <= 16'd963;
          lut[15240] <= 16'd1100;
          lut[15241] <= 16'd1237;
          lut[15242] <= 16'd1374;
          lut[15243] <= 16'd1510;
          lut[15244] <= 16'd1647;
          lut[15245] <= 16'd1783;
          lut[15246] <= 16'd1919;
          lut[15247] <= 16'd2054;
          lut[15248] <= 16'd2190;
          lut[15249] <= 16'd2325;
          lut[15250] <= 16'd2460;
          lut[15251] <= 16'd2594;
          lut[15252] <= 16'd2728;
          lut[15253] <= 16'd2862;
          lut[15254] <= 16'd2995;
          lut[15255] <= 16'd3128;
          lut[15256] <= 16'd3261;
          lut[15257] <= 16'd3393;
          lut[15258] <= 16'd3524;
          lut[15259] <= 16'd3655;
          lut[15260] <= 16'd3786;
          lut[15261] <= 16'd3916;
          lut[15262] <= 16'd4046;
          lut[15263] <= 16'd4175;
          lut[15264] <= 16'd4304;
          lut[15265] <= 16'd4432;
          lut[15266] <= 16'd4560;
          lut[15267] <= 16'd4687;
          lut[15268] <= 16'd4813;
          lut[15269] <= 16'd4939;
          lut[15270] <= 16'd5064;
          lut[15271] <= 16'd5189;
          lut[15272] <= 16'd5313;
          lut[15273] <= 16'd5436;
          lut[15274] <= 16'd5559;
          lut[15275] <= 16'd5681;
          lut[15276] <= 16'd5803;
          lut[15277] <= 16'd5923;
          lut[15278] <= 16'd6043;
          lut[15279] <= 16'd6163;
          lut[15280] <= 16'd6282;
          lut[15281] <= 16'd6400;
          lut[15282] <= 16'd6517;
          lut[15283] <= 16'd6634;
          lut[15284] <= 16'd6750;
          lut[15285] <= 16'd6865;
          lut[15286] <= 16'd6979;
          lut[15287] <= 16'd7093;
          lut[15288] <= 16'd7206;
          lut[15289] <= 16'd7319;
          lut[15290] <= 16'd7430;
          lut[15291] <= 16'd7541;
          lut[15292] <= 16'd7651;
          lut[15293] <= 16'd7761;
          lut[15294] <= 16'd7869;
          lut[15295] <= 16'd7977;
          lut[15296] <= 16'd8085;
          lut[15297] <= 16'd8191;
          lut[15298] <= 16'd8297;
          lut[15299] <= 16'd8402;
          lut[15300] <= 16'd8506;
          lut[15301] <= 16'd8609;
          lut[15302] <= 16'd8712;
          lut[15303] <= 16'd8814;
          lut[15304] <= 16'd8915;
          lut[15305] <= 16'd9015;
          lut[15306] <= 16'd9115;
          lut[15307] <= 16'd9214;
          lut[15308] <= 16'd9312;
          lut[15309] <= 16'd9409;
          lut[15310] <= 16'd9506;
          lut[15311] <= 16'd9602;
          lut[15312] <= 16'd9697;
          lut[15313] <= 16'd9792;
          lut[15314] <= 16'd9885;
          lut[15315] <= 16'd9978;
          lut[15316] <= 16'd10071;
          lut[15317] <= 16'd10162;
          lut[15318] <= 16'd10253;
          lut[15319] <= 16'd10343;
          lut[15320] <= 16'd10432;
          lut[15321] <= 16'd10521;
          lut[15322] <= 16'd10609;
          lut[15323] <= 16'd10696;
          lut[15324] <= 16'd10783;
          lut[15325] <= 16'd10869;
          lut[15326] <= 16'd10954;
          lut[15327] <= 16'd11038;
          lut[15328] <= 16'd11122;
          lut[15329] <= 16'd11205;
          lut[15330] <= 16'd11287;
          lut[15331] <= 16'd11369;
          lut[15332] <= 16'd11450;
          lut[15333] <= 16'd11530;
          lut[15334] <= 16'd11610;
          lut[15335] <= 16'd11689;
          lut[15336] <= 16'd11768;
          lut[15337] <= 16'd11845;
          lut[15338] <= 16'd11922;
          lut[15339] <= 16'd11999;
          lut[15340] <= 16'd12075;
          lut[15341] <= 16'd12150;
          lut[15342] <= 16'd12224;
          lut[15343] <= 16'd12298;
          lut[15344] <= 16'd12372;
          lut[15345] <= 16'd12444;
          lut[15346] <= 16'd12516;
          lut[15347] <= 16'd12588;
          lut[15348] <= 16'd12659;
          lut[15349] <= 16'd12729;
          lut[15350] <= 16'd12799;
          lut[15351] <= 16'd12868;
          lut[15352] <= 16'd12937;
          lut[15353] <= 16'd13004;
          lut[15354] <= 16'd13072;
          lut[15355] <= 16'd13139;
          lut[15356] <= 16'd13205;
          lut[15357] <= 16'd13271;
          lut[15358] <= 16'd13336;
          lut[15359] <= 16'd13401;
          lut[15360] <= 0;
          lut[15361] <= 16'd137;
          lut[15362] <= 16'd273;
          lut[15363] <= 16'd410;
          lut[15364] <= 16'd546;
          lut[15365] <= 16'd682;
          lut[15366] <= 16'd819;
          lut[15367] <= 16'd955;
          lut[15368] <= 16'd1091;
          lut[15369] <= 16'd1227;
          lut[15370] <= 16'd1362;
          lut[15371] <= 16'd1498;
          lut[15372] <= 16'd1633;
          lut[15373] <= 16'd1768;
          lut[15374] <= 16'd1903;
          lut[15375] <= 16'd2037;
          lut[15376] <= 16'd2172;
          lut[15377] <= 16'd2306;
          lut[15378] <= 16'd2439;
          lut[15379] <= 16'd2573;
          lut[15380] <= 16'd2706;
          lut[15381] <= 16'd2838;
          lut[15382] <= 16'd2971;
          lut[15383] <= 16'd3103;
          lut[15384] <= 16'd3234;
          lut[15385] <= 16'd3365;
          lut[15386] <= 16'd3496;
          lut[15387] <= 16'd3626;
          lut[15388] <= 16'd3756;
          lut[15389] <= 16'd3885;
          lut[15390] <= 16'd4014;
          lut[15391] <= 16'd4142;
          lut[15392] <= 16'd4270;
          lut[15393] <= 16'd4397;
          lut[15394] <= 16'd4524;
          lut[15395] <= 16'd4650;
          lut[15396] <= 16'd4775;
          lut[15397] <= 16'd4900;
          lut[15398] <= 16'd5025;
          lut[15399] <= 16'd5148;
          lut[15400] <= 16'd5272;
          lut[15401] <= 16'd5394;
          lut[15402] <= 16'd5516;
          lut[15403] <= 16'd5637;
          lut[15404] <= 16'd5758;
          lut[15405] <= 16'd5878;
          lut[15406] <= 16'd5997;
          lut[15407] <= 16'd6116;
          lut[15408] <= 16'd6234;
          lut[15409] <= 16'd6352;
          lut[15410] <= 16'd6468;
          lut[15411] <= 16'd6584;
          lut[15412] <= 16'd6700;
          lut[15413] <= 16'd6814;
          lut[15414] <= 16'd6928;
          lut[15415] <= 16'd7041;
          lut[15416] <= 16'd7154;
          lut[15417] <= 16'd7265;
          lut[15418] <= 16'd7376;
          lut[15419] <= 16'd7487;
          lut[15420] <= 16'd7596;
          lut[15421] <= 16'd7705;
          lut[15422] <= 16'd7813;
          lut[15423] <= 16'd7921;
          lut[15424] <= 16'd8027;
          lut[15425] <= 16'd8133;
          lut[15426] <= 16'd8239;
          lut[15427] <= 16'd8343;
          lut[15428] <= 16'd8447;
          lut[15429] <= 16'd8550;
          lut[15430] <= 16'd8652;
          lut[15431] <= 16'd8753;
          lut[15432] <= 16'd8854;
          lut[15433] <= 16'd8954;
          lut[15434] <= 16'd9054;
          lut[15435] <= 16'd9152;
          lut[15436] <= 16'd9250;
          lut[15437] <= 16'd9347;
          lut[15438] <= 16'd9443;
          lut[15439] <= 16'd9539;
          lut[15440] <= 16'd9634;
          lut[15441] <= 16'd9728;
          lut[15442] <= 16'd9821;
          lut[15443] <= 16'd9914;
          lut[15444] <= 16'd10006;
          lut[15445] <= 16'd10097;
          lut[15446] <= 16'd10188;
          lut[15447] <= 16'd10278;
          lut[15448] <= 16'd10367;
          lut[15449] <= 16'd10455;
          lut[15450] <= 16'd10543;
          lut[15451] <= 16'd10630;
          lut[15452] <= 16'd10716;
          lut[15453] <= 16'd10802;
          lut[15454] <= 16'd10887;
          lut[15455] <= 16'd10971;
          lut[15456] <= 16'd11055;
          lut[15457] <= 16'd11138;
          lut[15458] <= 16'd11220;
          lut[15459] <= 16'd11302;
          lut[15460] <= 16'd11383;
          lut[15461] <= 16'd11463;
          lut[15462] <= 16'd11542;
          lut[15463] <= 16'd11621;
          lut[15464] <= 16'd11700;
          lut[15465] <= 16'd11777;
          lut[15466] <= 16'd11854;
          lut[15467] <= 16'd11931;
          lut[15468] <= 16'd12006;
          lut[15469] <= 16'd12082;
          lut[15470] <= 16'd12156;
          lut[15471] <= 16'd12230;
          lut[15472] <= 16'd12303;
          lut[15473] <= 16'd12376;
          lut[15474] <= 16'd12448;
          lut[15475] <= 16'd12519;
          lut[15476] <= 16'd12590;
          lut[15477] <= 16'd12661;
          lut[15478] <= 16'd12730;
          lut[15479] <= 16'd12799;
          lut[15480] <= 16'd12868;
          lut[15481] <= 16'd12936;
          lut[15482] <= 16'd13003;
          lut[15483] <= 16'd13070;
          lut[15484] <= 16'd13137;
          lut[15485] <= 16'd13202;
          lut[15486] <= 16'd13267;
          lut[15487] <= 16'd13332;
          lut[15488] <= 0;
          lut[15489] <= 16'd135;
          lut[15490] <= 16'd271;
          lut[15491] <= 16'd406;
          lut[15492] <= 16'd541;
          lut[15493] <= 16'd677;
          lut[15494] <= 16'd812;
          lut[15495] <= 16'd947;
          lut[15496] <= 16'd1082;
          lut[15497] <= 16'd1216;
          lut[15498] <= 16'd1351;
          lut[15499] <= 16'd1485;
          lut[15500] <= 16'd1620;
          lut[15501] <= 16'd1754;
          lut[15502] <= 16'd1887;
          lut[15503] <= 16'd2021;
          lut[15504] <= 16'd2154;
          lut[15505] <= 16'd2287;
          lut[15506] <= 16'd2420;
          lut[15507] <= 16'd2552;
          lut[15508] <= 16'd2684;
          lut[15509] <= 16'd2815;
          lut[15510] <= 16'd2947;
          lut[15511] <= 16'd3078;
          lut[15512] <= 16'd3208;
          lut[15513] <= 16'd3338;
          lut[15514] <= 16'd3468;
          lut[15515] <= 16'd3597;
          lut[15516] <= 16'd3726;
          lut[15517] <= 16'd3854;
          lut[15518] <= 16'd3982;
          lut[15519] <= 16'd4109;
          lut[15520] <= 16'd4236;
          lut[15521] <= 16'd4362;
          lut[15522] <= 16'd4488;
          lut[15523] <= 16'd4613;
          lut[15524] <= 16'd4738;
          lut[15525] <= 16'd4862;
          lut[15526] <= 16'd4986;
          lut[15527] <= 16'd5109;
          lut[15528] <= 16'd5231;
          lut[15529] <= 16'd5353;
          lut[15530] <= 16'd5474;
          lut[15531] <= 16'd5594;
          lut[15532] <= 16'd5714;
          lut[15533] <= 16'd5834;
          lut[15534] <= 16'd5952;
          lut[15535] <= 16'd6070;
          lut[15536] <= 16'd6187;
          lut[15537] <= 16'd6304;
          lut[15538] <= 16'd6420;
          lut[15539] <= 16'd6535;
          lut[15540] <= 16'd6650;
          lut[15541] <= 16'd6764;
          lut[15542] <= 16'd6877;
          lut[15543] <= 16'd6990;
          lut[15544] <= 16'd7102;
          lut[15545] <= 16'd7213;
          lut[15546] <= 16'd7323;
          lut[15547] <= 16'd7433;
          lut[15548] <= 16'd7542;
          lut[15549] <= 16'd7650;
          lut[15550] <= 16'd7758;
          lut[15551] <= 16'd7865;
          lut[15552] <= 16'd7971;
          lut[15553] <= 16'd8077;
          lut[15554] <= 16'd8181;
          lut[15555] <= 16'd8285;
          lut[15556] <= 16'd8389;
          lut[15557] <= 16'd8491;
          lut[15558] <= 16'd8593;
          lut[15559] <= 16'd8694;
          lut[15560] <= 16'd8794;
          lut[15561] <= 16'd8894;
          lut[15562] <= 16'd8993;
          lut[15563] <= 16'd9091;
          lut[15564] <= 16'd9189;
          lut[15565] <= 16'd9285;
          lut[15566] <= 16'd9381;
          lut[15567] <= 16'd9477;
          lut[15568] <= 16'd9571;
          lut[15569] <= 16'd9665;
          lut[15570] <= 16'd9758;
          lut[15571] <= 16'd9851;
          lut[15572] <= 16'd9942;
          lut[15573] <= 16'd10033;
          lut[15574] <= 16'd10124;
          lut[15575] <= 16'd10213;
          lut[15576] <= 16'd10302;
          lut[15577] <= 16'd10390;
          lut[15578] <= 16'd10478;
          lut[15579] <= 16'd10565;
          lut[15580] <= 16'd10651;
          lut[15581] <= 16'd10736;
          lut[15582] <= 16'd10821;
          lut[15583] <= 16'd10905;
          lut[15584] <= 16'd10989;
          lut[15585] <= 16'd11071;
          lut[15586] <= 16'd11154;
          lut[15587] <= 16'd11235;
          lut[15588] <= 16'd11316;
          lut[15589] <= 16'd11396;
          lut[15590] <= 16'd11475;
          lut[15591] <= 16'd11554;
          lut[15592] <= 16'd11632;
          lut[15593] <= 16'd11710;
          lut[15594] <= 16'd11787;
          lut[15595] <= 16'd11863;
          lut[15596] <= 16'd11939;
          lut[15597] <= 16'd12014;
          lut[15598] <= 16'd12088;
          lut[15599] <= 16'd12162;
          lut[15600] <= 16'd12235;
          lut[15601] <= 16'd12308;
          lut[15602] <= 16'd12380;
          lut[15603] <= 16'd12452;
          lut[15604] <= 16'd12522;
          lut[15605] <= 16'd12593;
          lut[15606] <= 16'd12662;
          lut[15607] <= 16'd12731;
          lut[15608] <= 16'd12800;
          lut[15609] <= 16'd12868;
          lut[15610] <= 16'd12935;
          lut[15611] <= 16'd13002;
          lut[15612] <= 16'd13069;
          lut[15613] <= 16'd13134;
          lut[15614] <= 16'd13200;
          lut[15615] <= 16'd13264;
          lut[15616] <= 0;
          lut[15617] <= 16'd134;
          lut[15618] <= 16'd269;
          lut[15619] <= 16'd403;
          lut[15620] <= 16'd537;
          lut[15621] <= 16'd671;
          lut[15622] <= 16'd805;
          lut[15623] <= 16'd939;
          lut[15624] <= 16'd1073;
          lut[15625] <= 16'd1206;
          lut[15626] <= 16'd1340;
          lut[15627] <= 16'd1473;
          lut[15628] <= 16'd1606;
          lut[15629] <= 16'd1739;
          lut[15630] <= 16'd1872;
          lut[15631] <= 16'd2004;
          lut[15632] <= 16'd2137;
          lut[15633] <= 16'd2268;
          lut[15634] <= 16'd2400;
          lut[15635] <= 16'd2531;
          lut[15636] <= 16'd2662;
          lut[15637] <= 16'd2793;
          lut[15638] <= 16'd2923;
          lut[15639] <= 16'd3053;
          lut[15640] <= 16'd3182;
          lut[15641] <= 16'd3312;
          lut[15642] <= 16'd3440;
          lut[15643] <= 16'd3568;
          lut[15644] <= 16'd3696;
          lut[15645] <= 16'd3824;
          lut[15646] <= 16'd3950;
          lut[15647] <= 16'd4077;
          lut[15648] <= 16'd4203;
          lut[15649] <= 16'd4328;
          lut[15650] <= 16'd4453;
          lut[15651] <= 16'd4577;
          lut[15652] <= 16'd4701;
          lut[15653] <= 16'd4824;
          lut[15654] <= 16'd4947;
          lut[15655] <= 16'd5069;
          lut[15656] <= 16'd5191;
          lut[15657] <= 16'd5312;
          lut[15658] <= 16'd5432;
          lut[15659] <= 16'd5552;
          lut[15660] <= 16'd5671;
          lut[15661] <= 16'd5790;
          lut[15662] <= 16'd5908;
          lut[15663] <= 16'd6025;
          lut[15664] <= 16'd6141;
          lut[15665] <= 16'd6257;
          lut[15666] <= 16'd6373;
          lut[15667] <= 16'd6487;
          lut[15668] <= 16'd6601;
          lut[15669] <= 16'd6715;
          lut[15670] <= 16'd6827;
          lut[15671] <= 16'd6939;
          lut[15672] <= 16'd7050;
          lut[15673] <= 16'd7161;
          lut[15674] <= 16'd7271;
          lut[15675] <= 16'd7380;
          lut[15676] <= 16'd7489;
          lut[15677] <= 16'd7596;
          lut[15678] <= 16'd7703;
          lut[15679] <= 16'd7810;
          lut[15680] <= 16'd7916;
          lut[15681] <= 16'd8020;
          lut[15682] <= 16'd8125;
          lut[15683] <= 16'd8228;
          lut[15684] <= 16'd8331;
          lut[15685] <= 16'd8433;
          lut[15686] <= 16'd8535;
          lut[15687] <= 16'd8635;
          lut[15688] <= 16'd8735;
          lut[15689] <= 16'd8834;
          lut[15690] <= 16'd8933;
          lut[15691] <= 16'd9031;
          lut[15692] <= 16'd9128;
          lut[15693] <= 16'd9224;
          lut[15694] <= 16'd9320;
          lut[15695] <= 16'd9415;
          lut[15696] <= 16'd9509;
          lut[15697] <= 16'd9603;
          lut[15698] <= 16'd9696;
          lut[15699] <= 16'd9788;
          lut[15700] <= 16'd9879;
          lut[15701] <= 16'd9970;
          lut[15702] <= 16'd10060;
          lut[15703] <= 16'd10149;
          lut[15704] <= 16'd10238;
          lut[15705] <= 16'd10326;
          lut[15706] <= 16'd10413;
          lut[15707] <= 16'd10500;
          lut[15708] <= 16'd10586;
          lut[15709] <= 16'd10671;
          lut[15710] <= 16'd10756;
          lut[15711] <= 16'd10840;
          lut[15712] <= 16'd10923;
          lut[15713] <= 16'd11006;
          lut[15714] <= 16'd11088;
          lut[15715] <= 16'd11169;
          lut[15716] <= 16'd11250;
          lut[15717] <= 16'd11330;
          lut[15718] <= 16'd11409;
          lut[15719] <= 16'd11488;
          lut[15720] <= 16'd11566;
          lut[15721] <= 16'd11643;
          lut[15722] <= 16'd11720;
          lut[15723] <= 16'd11796;
          lut[15724] <= 16'd11872;
          lut[15725] <= 16'd11947;
          lut[15726] <= 16'd12021;
          lut[15727] <= 16'd12095;
          lut[15728] <= 16'd12168;
          lut[15729] <= 16'd12241;
          lut[15730] <= 16'd12313;
          lut[15731] <= 16'd12384;
          lut[15732] <= 16'd12455;
          lut[15733] <= 16'd12525;
          lut[15734] <= 16'd12595;
          lut[15735] <= 16'd12664;
          lut[15736] <= 16'd12733;
          lut[15737] <= 16'd12801;
          lut[15738] <= 16'd12868;
          lut[15739] <= 16'd12935;
          lut[15740] <= 16'd13001;
          lut[15741] <= 16'd13067;
          lut[15742] <= 16'd13132;
          lut[15743] <= 16'd13197;
          lut[15744] <= 0;
          lut[15745] <= 16'd133;
          lut[15746] <= 16'd266;
          lut[15747] <= 16'd400;
          lut[15748] <= 16'd533;
          lut[15749] <= 16'd666;
          lut[15750] <= 16'd799;
          lut[15751] <= 16'd931;
          lut[15752] <= 16'd1064;
          lut[15753] <= 16'd1197;
          lut[15754] <= 16'd1329;
          lut[15755] <= 16'd1461;
          lut[15756] <= 16'd1593;
          lut[15757] <= 16'd1725;
          lut[15758] <= 16'd1857;
          lut[15759] <= 16'd1988;
          lut[15760] <= 16'd2119;
          lut[15761] <= 16'd2250;
          lut[15762] <= 16'd2381;
          lut[15763] <= 16'd2511;
          lut[15764] <= 16'd2641;
          lut[15765] <= 16'd2771;
          lut[15766] <= 16'd2900;
          lut[15767] <= 16'd3029;
          lut[15768] <= 16'd3157;
          lut[15769] <= 16'd3285;
          lut[15770] <= 16'd3413;
          lut[15771] <= 16'd3540;
          lut[15772] <= 16'd3667;
          lut[15773] <= 16'd3794;
          lut[15774] <= 16'd3920;
          lut[15775] <= 16'd4045;
          lut[15776] <= 16'd4170;
          lut[15777] <= 16'd4295;
          lut[15778] <= 16'd4419;
          lut[15779] <= 16'd4542;
          lut[15780] <= 16'd4665;
          lut[15781] <= 16'd4787;
          lut[15782] <= 16'd4909;
          lut[15783] <= 16'd5031;
          lut[15784] <= 16'd5151;
          lut[15785] <= 16'd5272;
          lut[15786] <= 16'd5391;
          lut[15787] <= 16'd5510;
          lut[15788] <= 16'd5629;
          lut[15789] <= 16'd5746;
          lut[15790] <= 16'd5863;
          lut[15791] <= 16'd5980;
          lut[15792] <= 16'd6096;
          lut[15793] <= 16'd6211;
          lut[15794] <= 16'd6326;
          lut[15795] <= 16'd6440;
          lut[15796] <= 16'd6553;
          lut[15797] <= 16'd6666;
          lut[15798] <= 16'd6778;
          lut[15799] <= 16'd6889;
          lut[15800] <= 16'd7000;
          lut[15801] <= 16'd7110;
          lut[15802] <= 16'd7219;
          lut[15803] <= 16'd7328;
          lut[15804] <= 16'd7436;
          lut[15805] <= 16'd7543;
          lut[15806] <= 16'd7650;
          lut[15807] <= 16'd7755;
          lut[15808] <= 16'd7861;
          lut[15809] <= 16'd7965;
          lut[15810] <= 16'd8069;
          lut[15811] <= 16'd8172;
          lut[15812] <= 16'd8274;
          lut[15813] <= 16'd8376;
          lut[15814] <= 16'd8477;
          lut[15815] <= 16'd8577;
          lut[15816] <= 16'd8677;
          lut[15817] <= 16'd8776;
          lut[15818] <= 16'd8874;
          lut[15819] <= 16'd8971;
          lut[15820] <= 16'd9068;
          lut[15821] <= 16'd9164;
          lut[15822] <= 16'd9259;
          lut[15823] <= 16'd9354;
          lut[15824] <= 16'd9448;
          lut[15825] <= 16'd9541;
          lut[15826] <= 16'd9634;
          lut[15827] <= 16'd9726;
          lut[15828] <= 16'd9817;
          lut[15829] <= 16'd9907;
          lut[15830] <= 16'd9997;
          lut[15831] <= 16'd10086;
          lut[15832] <= 16'd10175;
          lut[15833] <= 16'd10263;
          lut[15834] <= 16'd10350;
          lut[15835] <= 16'd10436;
          lut[15836] <= 16'd10522;
          lut[15837] <= 16'd10607;
          lut[15838] <= 16'd10691;
          lut[15839] <= 16'd10775;
          lut[15840] <= 16'd10858;
          lut[15841] <= 16'd10941;
          lut[15842] <= 16'd11022;
          lut[15843] <= 16'd11104;
          lut[15844] <= 16'd11184;
          lut[15845] <= 16'd11264;
          lut[15846] <= 16'd11343;
          lut[15847] <= 16'd11422;
          lut[15848] <= 16'd11500;
          lut[15849] <= 16'd11577;
          lut[15850] <= 16'd11654;
          lut[15851] <= 16'd11730;
          lut[15852] <= 16'd11806;
          lut[15853] <= 16'd11880;
          lut[15854] <= 16'd11955;
          lut[15855] <= 16'd12028;
          lut[15856] <= 16'd12102;
          lut[15857] <= 16'd12174;
          lut[15858] <= 16'd12246;
          lut[15859] <= 16'd12317;
          lut[15860] <= 16'd12388;
          lut[15861] <= 16'd12458;
          lut[15862] <= 16'd12528;
          lut[15863] <= 16'd12597;
          lut[15864] <= 16'd12666;
          lut[15865] <= 16'd12734;
          lut[15866] <= 16'd12801;
          lut[15867] <= 16'd12868;
          lut[15868] <= 16'd12934;
          lut[15869] <= 16'd13000;
          lut[15870] <= 16'd13065;
          lut[15871] <= 16'd13130;
          lut[15872] <= 0;
          lut[15873] <= 16'd132;
          lut[15874] <= 16'd264;
          lut[15875] <= 16'd396;
          lut[15876] <= 16'd528;
          lut[15877] <= 16'd660;
          lut[15878] <= 16'd792;
          lut[15879] <= 16'd924;
          lut[15880] <= 16'd1056;
          lut[15881] <= 16'd1187;
          lut[15882] <= 16'd1318;
          lut[15883] <= 16'd1450;
          lut[15884] <= 16'd1581;
          lut[15885] <= 16'd1711;
          lut[15886] <= 16'd1842;
          lut[15887] <= 16'd1972;
          lut[15888] <= 16'd2102;
          lut[15889] <= 16'd2232;
          lut[15890] <= 16'd2362;
          lut[15891] <= 16'd2491;
          lut[15892] <= 16'd2620;
          lut[15893] <= 16'd2749;
          lut[15894] <= 16'd2877;
          lut[15895] <= 16'd3005;
          lut[15896] <= 16'd3132;
          lut[15897] <= 16'd3260;
          lut[15898] <= 16'd3386;
          lut[15899] <= 16'd3513;
          lut[15900] <= 16'd3639;
          lut[15901] <= 16'd3764;
          lut[15902] <= 16'd3889;
          lut[15903] <= 16'd4014;
          lut[15904] <= 16'd4138;
          lut[15905] <= 16'd4261;
          lut[15906] <= 16'd4385;
          lut[15907] <= 16'd4507;
          lut[15908] <= 16'd4629;
          lut[15909] <= 16'd4751;
          lut[15910] <= 16'd4872;
          lut[15911] <= 16'd4993;
          lut[15912] <= 16'd5112;
          lut[15913] <= 16'd5232;
          lut[15914] <= 16'd5351;
          lut[15915] <= 16'd5469;
          lut[15916] <= 16'd5587;
          lut[15917] <= 16'd5704;
          lut[15918] <= 16'd5820;
          lut[15919] <= 16'd5936;
          lut[15920] <= 16'd6051;
          lut[15921] <= 16'd6166;
          lut[15922] <= 16'd6280;
          lut[15923] <= 16'd6393;
          lut[15924] <= 16'd6506;
          lut[15925] <= 16'd6618;
          lut[15926] <= 16'd6729;
          lut[15927] <= 16'd6840;
          lut[15928] <= 16'd6950;
          lut[15929] <= 16'd7059;
          lut[15930] <= 16'd7168;
          lut[15931] <= 16'd7276;
          lut[15932] <= 16'd7384;
          lut[15933] <= 16'd7490;
          lut[15934] <= 16'd7596;
          lut[15935] <= 16'd7702;
          lut[15936] <= 16'd7806;
          lut[15937] <= 16'd7910;
          lut[15938] <= 16'd8014;
          lut[15939] <= 16'd8116;
          lut[15940] <= 16'd8218;
          lut[15941] <= 16'd8320;
          lut[15942] <= 16'd8420;
          lut[15943] <= 16'd8520;
          lut[15944] <= 16'd8619;
          lut[15945] <= 16'd8718;
          lut[15946] <= 16'd8815;
          lut[15947] <= 16'd8912;
          lut[15948] <= 16'd9009;
          lut[15949] <= 16'd9104;
          lut[15950] <= 16'd9200;
          lut[15951] <= 16'd9294;
          lut[15952] <= 16'd9387;
          lut[15953] <= 16'd9480;
          lut[15954] <= 16'd9573;
          lut[15955] <= 16'd9664;
          lut[15956] <= 16'd9755;
          lut[15957] <= 16'd9845;
          lut[15958] <= 16'd9935;
          lut[15959] <= 16'd10024;
          lut[15960] <= 16'd10112;
          lut[15961] <= 16'd10200;
          lut[15962] <= 16'd10286;
          lut[15963] <= 16'd10373;
          lut[15964] <= 16'd10458;
          lut[15965] <= 16'd10543;
          lut[15966] <= 16'd10627;
          lut[15967] <= 16'd10711;
          lut[15968] <= 16'd10794;
          lut[15969] <= 16'd10876;
          lut[15970] <= 16'd10958;
          lut[15971] <= 16'd11039;
          lut[15972] <= 16'd11119;
          lut[15973] <= 16'd11199;
          lut[15974] <= 16'd11278;
          lut[15975] <= 16'd11357;
          lut[15976] <= 16'd11434;
          lut[15977] <= 16'd11512;
          lut[15978] <= 16'd11588;
          lut[15979] <= 16'd11664;
          lut[15980] <= 16'd11740;
          lut[15981] <= 16'd11815;
          lut[15982] <= 16'd11889;
          lut[15983] <= 16'd11963;
          lut[15984] <= 16'd12036;
          lut[15985] <= 16'd12108;
          lut[15986] <= 16'd12180;
          lut[15987] <= 16'd12251;
          lut[15988] <= 16'd12322;
          lut[15989] <= 16'd12392;
          lut[15990] <= 16'd12462;
          lut[15991] <= 16'd12531;
          lut[15992] <= 16'd12599;
          lut[15993] <= 16'd12667;
          lut[15994] <= 16'd12735;
          lut[15995] <= 16'd12802;
          lut[15996] <= 16'd12868;
          lut[15997] <= 16'd12934;
          lut[15998] <= 16'd12999;
          lut[15999] <= 16'd13064;
          lut[16000] <= 0;
          lut[16001] <= 16'd131;
          lut[16002] <= 16'd262;
          lut[16003] <= 16'd393;
          lut[16004] <= 16'd524;
          lut[16005] <= 16'd655;
          lut[16006] <= 16'd786;
          lut[16007] <= 16'd917;
          lut[16008] <= 16'd1047;
          lut[16009] <= 16'd1178;
          lut[16010] <= 16'd1308;
          lut[16011] <= 16'd1438;
          lut[16012] <= 16'd1568;
          lut[16013] <= 16'd1698;
          lut[16014] <= 16'd1827;
          lut[16015] <= 16'd1957;
          lut[16016] <= 16'd2086;
          lut[16017] <= 16'd2215;
          lut[16018] <= 16'd2343;
          lut[16019] <= 16'd2471;
          lut[16020] <= 16'd2599;
          lut[16021] <= 16'd2727;
          lut[16022] <= 16'd2854;
          lut[16023] <= 16'd2981;
          lut[16024] <= 16'd3108;
          lut[16025] <= 16'd3234;
          lut[16026] <= 16'd3360;
          lut[16027] <= 16'd3485;
          lut[16028] <= 16'd3610;
          lut[16029] <= 16'd3735;
          lut[16030] <= 16'd3859;
          lut[16031] <= 16'd3983;
          lut[16032] <= 16'd4106;
          lut[16033] <= 16'd4229;
          lut[16034] <= 16'd4351;
          lut[16035] <= 16'd4473;
          lut[16036] <= 16'd4594;
          lut[16037] <= 16'd4715;
          lut[16038] <= 16'd4835;
          lut[16039] <= 16'd4955;
          lut[16040] <= 16'd5074;
          lut[16041] <= 16'd5193;
          lut[16042] <= 16'd5311;
          lut[16043] <= 16'd5428;
          lut[16044] <= 16'd5545;
          lut[16045] <= 16'd5662;
          lut[16046] <= 16'd5777;
          lut[16047] <= 16'd5892;
          lut[16048] <= 16'd6007;
          lut[16049] <= 16'd6121;
          lut[16050] <= 16'd6234;
          lut[16051] <= 16'd6347;
          lut[16052] <= 16'd6459;
          lut[16053] <= 16'd6570;
          lut[16054] <= 16'd6681;
          lut[16055] <= 16'd6791;
          lut[16056] <= 16'd6901;
          lut[16057] <= 16'd7010;
          lut[16058] <= 16'd7118;
          lut[16059] <= 16'd7225;
          lut[16060] <= 16'd7332;
          lut[16061] <= 16'd7438;
          lut[16062] <= 16'd7544;
          lut[16063] <= 16'd7649;
          lut[16064] <= 16'd7753;
          lut[16065] <= 16'd7856;
          lut[16066] <= 16'd7959;
          lut[16067] <= 16'd8061;
          lut[16068] <= 16'd8163;
          lut[16069] <= 16'd8264;
          lut[16070] <= 16'd8364;
          lut[16071] <= 16'd8463;
          lut[16072] <= 16'd8562;
          lut[16073] <= 16'd8660;
          lut[16074] <= 16'd8758;
          lut[16075] <= 16'd8854;
          lut[16076] <= 16'd8950;
          lut[16077] <= 16'd9046;
          lut[16078] <= 16'd9140;
          lut[16079] <= 16'd9234;
          lut[16080] <= 16'd9328;
          lut[16081] <= 16'd9420;
          lut[16082] <= 16'd9512;
          lut[16083] <= 16'd9604;
          lut[16084] <= 16'd9694;
          lut[16085] <= 16'd9784;
          lut[16086] <= 16'd9873;
          lut[16087] <= 16'd9962;
          lut[16088] <= 16'd10050;
          lut[16089] <= 16'd10137;
          lut[16090] <= 16'd10224;
          lut[16091] <= 16'd10310;
          lut[16092] <= 16'd10395;
          lut[16093] <= 16'd10480;
          lut[16094] <= 16'd10564;
          lut[16095] <= 16'd10647;
          lut[16096] <= 16'd10730;
          lut[16097] <= 16'd10812;
          lut[16098] <= 16'd10894;
          lut[16099] <= 16'd10975;
          lut[16100] <= 16'd11055;
          lut[16101] <= 16'd11135;
          lut[16102] <= 16'd11214;
          lut[16103] <= 16'd11292;
          lut[16104] <= 16'd11370;
          lut[16105] <= 16'd11447;
          lut[16106] <= 16'd11523;
          lut[16107] <= 16'd11599;
          lut[16108] <= 16'd11675;
          lut[16109] <= 16'd11749;
          lut[16110] <= 16'd11824;
          lut[16111] <= 16'd11897;
          lut[16112] <= 16'd11970;
          lut[16113] <= 16'd12043;
          lut[16114] <= 16'd12114;
          lut[16115] <= 16'd12186;
          lut[16116] <= 16'd12256;
          lut[16117] <= 16'd12327;
          lut[16118] <= 16'd12396;
          lut[16119] <= 16'd12465;
          lut[16120] <= 16'd12534;
          lut[16121] <= 16'd12602;
          lut[16122] <= 16'd12669;
          lut[16123] <= 16'd12736;
          lut[16124] <= 16'd12802;
          lut[16125] <= 16'd12868;
          lut[16126] <= 16'd12933;
          lut[16127] <= 16'd12998;
          lut[16128] <= 0;
          lut[16129] <= 16'd130;
          lut[16130] <= 16'd260;
          lut[16131] <= 16'd390;
          lut[16132] <= 16'd520;
          lut[16133] <= 16'd650;
          lut[16134] <= 16'd780;
          lut[16135] <= 16'd909;
          lut[16136] <= 16'd1039;
          lut[16137] <= 16'd1168;
          lut[16138] <= 16'd1298;
          lut[16139] <= 16'd1427;
          lut[16140] <= 16'd1556;
          lut[16141] <= 16'd1684;
          lut[16142] <= 16'd1813;
          lut[16143] <= 16'd1941;
          lut[16144] <= 16'd2069;
          lut[16145] <= 16'd2197;
          lut[16146] <= 16'd2325;
          lut[16147] <= 16'd2452;
          lut[16148] <= 16'd2579;
          lut[16149] <= 16'd2706;
          lut[16150] <= 16'd2832;
          lut[16151] <= 16'd2958;
          lut[16152] <= 16'd3084;
          lut[16153] <= 16'd3209;
          lut[16154] <= 16'd3334;
          lut[16155] <= 16'd3459;
          lut[16156] <= 16'd3583;
          lut[16157] <= 16'd3706;
          lut[16158] <= 16'd3830;
          lut[16159] <= 16'd3952;
          lut[16160] <= 16'd4075;
          lut[16161] <= 16'd4197;
          lut[16162] <= 16'd4318;
          lut[16163] <= 16'd4439;
          lut[16164] <= 16'd4560;
          lut[16165] <= 16'd4680;
          lut[16166] <= 16'd4799;
          lut[16167] <= 16'd4918;
          lut[16168] <= 16'd5036;
          lut[16169] <= 16'd5154;
          lut[16170] <= 16'd5272;
          lut[16171] <= 16'd5388;
          lut[16172] <= 16'd5504;
          lut[16173] <= 16'd5620;
          lut[16174] <= 16'd5735;
          lut[16175] <= 16'd5850;
          lut[16176] <= 16'd5963;
          lut[16177] <= 16'd6077;
          lut[16178] <= 16'd6189;
          lut[16179] <= 16'd6301;
          lut[16180] <= 16'd6413;
          lut[16181] <= 16'd6524;
          lut[16182] <= 16'd6634;
          lut[16183] <= 16'd6743;
          lut[16184] <= 16'd6852;
          lut[16185] <= 16'd6960;
          lut[16186] <= 16'd7068;
          lut[16187] <= 16'd7175;
          lut[16188] <= 16'd7281;
          lut[16189] <= 16'd7387;
          lut[16190] <= 16'd7492;
          lut[16191] <= 16'd7596;
          lut[16192] <= 16'd7700;
          lut[16193] <= 16'd7803;
          lut[16194] <= 16'd7905;
          lut[16195] <= 16'd8007;
          lut[16196] <= 16'd8108;
          lut[16197] <= 16'd8209;
          lut[16198] <= 16'd8308;
          lut[16199] <= 16'd8407;
          lut[16200] <= 16'd8506;
          lut[16201] <= 16'd8603;
          lut[16202] <= 16'd8700;
          lut[16203] <= 16'd8797;
          lut[16204] <= 16'd8892;
          lut[16205] <= 16'd8987;
          lut[16206] <= 16'd9082;
          lut[16207] <= 16'd9175;
          lut[16208] <= 16'd9268;
          lut[16209] <= 16'd9361;
          lut[16210] <= 16'd9452;
          lut[16211] <= 16'd9543;
          lut[16212] <= 16'd9634;
          lut[16213] <= 16'd9724;
          lut[16214] <= 16'd9813;
          lut[16215] <= 16'd9901;
          lut[16216] <= 16'd9989;
          lut[16217] <= 16'd10076;
          lut[16218] <= 16'd10162;
          lut[16219] <= 16'd10248;
          lut[16220] <= 16'd10333;
          lut[16221] <= 16'd10418;
          lut[16222] <= 16'd10501;
          lut[16223] <= 16'd10585;
          lut[16224] <= 16'd10667;
          lut[16225] <= 16'd10749;
          lut[16226] <= 16'd10831;
          lut[16227] <= 16'd10911;
          lut[16228] <= 16'd10991;
          lut[16229] <= 16'd11071;
          lut[16230] <= 16'd11150;
          lut[16231] <= 16'd11228;
          lut[16232] <= 16'd11306;
          lut[16233] <= 16'd11383;
          lut[16234] <= 16'd11459;
          lut[16235] <= 16'd11535;
          lut[16236] <= 16'd11610;
          lut[16237] <= 16'd11685;
          lut[16238] <= 16'd11759;
          lut[16239] <= 16'd11832;
          lut[16240] <= 16'd11905;
          lut[16241] <= 16'd11978;
          lut[16242] <= 16'd12049;
          lut[16243] <= 16'd12121;
          lut[16244] <= 16'd12191;
          lut[16245] <= 16'd12261;
          lut[16246] <= 16'd12331;
          lut[16247] <= 16'd12400;
          lut[16248] <= 16'd12468;
          lut[16249] <= 16'd12536;
          lut[16250] <= 16'd12604;
          lut[16251] <= 16'd12671;
          lut[16252] <= 16'd12737;
          lut[16253] <= 16'd12803;
          lut[16254] <= 16'd12868;
          lut[16255] <= 16'd12933;
          lut[16256] <= 0;
          lut[16257] <= 16'd129;
          lut[16258] <= 16'd258;
          lut[16259] <= 16'd387;
          lut[16260] <= 16'd516;
          lut[16261] <= 16'd645;
          lut[16262] <= 16'd773;
          lut[16263] <= 16'd902;
          lut[16264] <= 16'd1031;
          lut[16265] <= 16'd1159;
          lut[16266] <= 16'd1287;
          lut[16267] <= 16'd1416;
          lut[16268] <= 16'd1544;
          lut[16269] <= 16'd1671;
          lut[16270] <= 16'd1799;
          lut[16271] <= 16'd1926;
          lut[16272] <= 16'd2053;
          lut[16273] <= 16'd2180;
          lut[16274] <= 16'd2307;
          lut[16275] <= 16'd2433;
          lut[16276] <= 16'd2559;
          lut[16277] <= 16'd2685;
          lut[16278] <= 16'd2810;
          lut[16279] <= 16'd2935;
          lut[16280] <= 16'd3060;
          lut[16281] <= 16'd3184;
          lut[16282] <= 16'd3308;
          lut[16283] <= 16'd3432;
          lut[16284] <= 16'd3555;
          lut[16285] <= 16'd3678;
          lut[16286] <= 16'd3801;
          lut[16287] <= 16'd3923;
          lut[16288] <= 16'd4044;
          lut[16289] <= 16'd4165;
          lut[16290] <= 16'd4286;
          lut[16291] <= 16'd4406;
          lut[16292] <= 16'd4526;
          lut[16293] <= 16'd4645;
          lut[16294] <= 16'd4763;
          lut[16295] <= 16'd4882;
          lut[16296] <= 16'd4999;
          lut[16297] <= 16'd5116;
          lut[16298] <= 16'd5233;
          lut[16299] <= 16'd5349;
          lut[16300] <= 16'd5464;
          lut[16301] <= 16'd5579;
          lut[16302] <= 16'd5694;
          lut[16303] <= 16'd5807;
          lut[16304] <= 16'd5920;
          lut[16305] <= 16'd6033;
          lut[16306] <= 16'd6145;
          lut[16307] <= 16'd6256;
          lut[16308] <= 16'd6367;
          lut[16309] <= 16'd6477;
          lut[16310] <= 16'd6587;
          lut[16311] <= 16'd6696;
          lut[16312] <= 16'd6804;
          lut[16313] <= 16'd6912;
          lut[16314] <= 16'd7019;
          lut[16315] <= 16'd7125;
          lut[16316] <= 16'd7231;
          lut[16317] <= 16'd7336;
          lut[16318] <= 16'd7441;
          lut[16319] <= 16'd7545;
          lut[16320] <= 16'd7648;
          lut[16321] <= 16'd7750;
          lut[16322] <= 16'd7852;
          lut[16323] <= 16'd7954;
          lut[16324] <= 16'd8054;
          lut[16325] <= 16'd8154;
          lut[16326] <= 16'd8253;
          lut[16327] <= 16'd8352;
          lut[16328] <= 16'd8450;
          lut[16329] <= 16'd8547;
          lut[16330] <= 16'd8644;
          lut[16331] <= 16'd8740;
          lut[16332] <= 16'd8835;
          lut[16333] <= 16'd8930;
          lut[16334] <= 16'd9024;
          lut[16335] <= 16'd9117;
          lut[16336] <= 16'd9210;
          lut[16337] <= 16'd9302;
          lut[16338] <= 16'd9393;
          lut[16339] <= 16'd9484;
          lut[16340] <= 16'd9574;
          lut[16341] <= 16'd9664;
          lut[16342] <= 16'd9752;
          lut[16343] <= 16'd9840;
          lut[16344] <= 16'd9928;
          lut[16345] <= 16'd10015;
          lut[16346] <= 16'd10101;
          lut[16347] <= 16'd10187;
          lut[16348] <= 16'd10271;
          lut[16349] <= 16'd10356;
          lut[16350] <= 16'd10439;
          lut[16351] <= 16'd10522;
          lut[16352] <= 16'd10605;
          lut[16353] <= 16'd10687;
          lut[16354] <= 16'd10768;
          lut[16355] <= 16'd10848;
          lut[16356] <= 16'd10928;
          lut[16357] <= 16'd11008;
          lut[16358] <= 16'd11086;
          lut[16359] <= 16'd11164;
          lut[16360] <= 16'd11242;
          lut[16361] <= 16'd11319;
          lut[16362] <= 16'd11395;
          lut[16363] <= 16'd11471;
          lut[16364] <= 16'd11546;
          lut[16365] <= 16'd11621;
          lut[16366] <= 16'd11695;
          lut[16367] <= 16'd11768;
          lut[16368] <= 16'd11841;
          lut[16369] <= 16'd11913;
          lut[16370] <= 16'd11985;
          lut[16371] <= 16'd12056;
          lut[16372] <= 16'd12127;
          lut[16373] <= 16'd12197;
          lut[16374] <= 16'd12266;
          lut[16375] <= 16'd12335;
          lut[16376] <= 16'd12404;
          lut[16377] <= 16'd12472;
          lut[16378] <= 16'd12539;
          lut[16379] <= 16'd12606;
          lut[16380] <= 16'd12672;
          lut[16381] <= 16'd12738;
          lut[16382] <= 16'd12803;
          lut[16383] <= 16'd12868;
       end
    end
endmodule
